/*
input logic clock_10_i,
input logic reset_i,
input logic locked_i,
output logic reset_effectivo_o,


output logic [15:0] led_o,
input logic [15:0] sw_i,
input logic [3:0] btn_i,
output logic [6:0] segmentos_o,
output logic [7:0] anodos_o,
output logic dp_o,

output logic [10:0] instr_addr_bus_o,
input logic [31:0] instr_bus_i,

output logic [31:0] address_ext_o,
input logic [31:0] ext_bus_data_i,
output logic [31:0] ext_bus_data_o,
output logic        ext_bus_we_o,

output logic [9:0] ram_address_bus_o,
output logic        ram_we_o,
output logic [31:0] ram_data_in_o,
input logic [31:0] ram_data_out_i
*/

module microcontrolador_syn(clock_10_i, reset_i, locked_i, reset_effectivo_o, led_o, sw_i, btn_i, segmentos_o, anodos_o, dp_o, instr_addr_bus_o, instr_bus_i, address_ext_o, ext_bus_data_i, ext_bus_data_o, ext_bus_we_o, ram_address_bus_o, ram_we_o, ram_data_in_o, ram_data_out_i);
  reg [4:0] nr00000;
  reg [4:0] nr00001;
  wire nw00000;
  wire nw00001;
  wire nw00002;
  wire nw00003;
  wire nw00004;
  wire nw00005;
  wire nw00006;
  wire nw00007;
  wire nw00008;
  wire nw00009;
  wire nw00010;
  wire nw00011;
  wire nw00012;
  wire nw00013;
  wire nw00014;
  wire nw00015;
  wire nw00016;
  wire nw00017;
  wire nw00018;
  wire nw00019;
  wire nw00020;
  wire nw00021;
  wire nw00022;
  wire nw00023;
  wire nw00024;
  wire nw00025;
  wire nw00026;
  wire nw00027;
  wire nw00028;
  wire nw00029;
  wire nw00030;
  wire nw00031;
  wire nw00032;
  wire nw00033;
  wire nw00034;
  wire nw00035;
  wire nw00036;
  wire nw00037;
  wire nw00038;
  wire nw00039;
  wire nw00040;
  wire nw00041;
  wire nw00042;
  wire nw00043;
  wire nw00044;
  wire nw00045;
  wire nw00046;
  wire nw00047;
  wire nw00048;
  wire nw00049;
  wire nw00050;
  wire nw00051;
  wire nw00052;
  wire nw00053;
  wire nw00054;
  wire nw00055;
  wire nw00056;
  wire nw00057;
  wire nw00058;
  wire nw00059;
  wire nw00060;
  wire nw00061;
  wire nw00062;
  wire nw00063;
  wire nw00064;
  wire nw00065;
  wire nw00066;
  wire nw00067;
  wire nw00068;
  wire nw00069;
  wire nw00070;
  wire nw00071;
  wire nw00072;
  wire nw00073;
  wire nw00074;
  wire nw00075;
  wire nw00076;
  wire nw00077;
  wire nw00078;
  wire nw00079;
  wire nw00080;
  wire nw00081;
  wire nw00082;
  wire nw00083;
  wire nw00084;
  wire nw00085;
  wire nw00086;
  wire nw00087;
  wire nw00088;
  wire nw00089;
  wire nw00090;
  wire nw00091;
  wire nw00092;
  wire nw00093;
  wire nw00094;
  wire nw00095;
  wire nw00096;
  wire nw00097;
  wire nw00098;
  wire nw00099;
  wire nw00100;
  wire nw00101;
  wire nw00102;
  wire nw00103;
  wire nw00104;
  wire nw00105;
  wire nw00106;
  wire nw00107;
  wire nw00108;
  wire nw00109;
  wire nw00110;
  wire nw00111;
  wire nw00112;
  wire nw00113;
  wire nw00114;
  wire nw00115;
  wire nw00116;
  wire nw00117;
  wire nw00118;
  wire nw00119;
  wire nw00120;
  wire nw00121;
  wire nw00122;
  wire nw00123;
  wire nw00124;
  wire nw00125;
  wire nw00126;
  wire nw00127;
  wire nw00128;
  wire nw00129;
  wire nw00130;
  wire nw00131;
  wire nw00132;
  wire nw00133;
  wire nw00134;
  wire nw00135;
  wire nw00136;
  wire nw00137;
  wire nw00138;
  wire nw00139;
  wire nw00140;
  wire nw00141;
  wire nw00142;
  wire nw00143;
  wire nw00144;
  wire nw00145;
  wire nw00146;
  wire nw00147;
  wire nw00148;
  wire nw00149;
  wire nw00150;
  wire nw00151;
  wire nw00152;
  wire nw00153;
  wire nw00154;
  wire nw00155;
  wire nw00156;
  wire nw00157;
  wire nw00158;
  wire nw00159;
  wire nw00160;
  wire nw00161;
  wire nw00162;
  wire nw00163;
  wire nw00164;
  wire nw00165;
  wire nw00166;
  wire nw00167;
  wire nw00168;
  wire nw00169;
  wire nw00170;
  wire nw00171;
  wire nw00172;
  wire nw00173;
  wire nw00174;
  wire nw00175;
  wire nw00176;
  wire nw00177;
  wire nw00178;
  wire nw00179;
  wire nw00180;
  wire nw00181;
  wire nw00182;
  wire nw00183;
  wire nw00184;
  wire nw00185;
  wire nw00186;
  wire nw00187;
  wire nw00188;
  wire nw00189;
  wire nw00190;
  wire nw00191;
  wire nw00192;
  wire nw00193;
  wire nw00194;
  wire nw00195;
  wire nw00196;
  wire nw00197;
  wire nw00198;
  wire nw00199;
  wire nw00200;
  wire nw00201;
  wire nw00202;
  wire nw00203;
  wire nw00204;
  wire nw00205;
  wire nw00206;
  wire nw00207;
  wire nw00208;
  wire nw00209;
  wire nw00210;
  wire nw00211;
  wire nw00212;
  wire nw00213;
  wire nw00214;
  wire nw00215;
  wire nw00216;
  wire nw00217;
  wire nw00218;
  wire nw00219;
  wire nw00220;
  wire nw00221;
  wire nw00222;
  wire nw00223;
  wire nw00224;
  wire nw00225;
  wire nw00226;
  wire nw00227;
  wire nw00228;
  wire nw00229;
  wire nw00230;
  wire nw00231;
  wire nw00232;
  wire nw00233;
  wire nw00234;
  wire nw00235;
  wire nw00236;
  wire nw00237;
  wire nw00238;
  wire nw00239;
  wire nw00240;
  wire nw00241;
  wire nw00242;
  wire nw00243;
  wire nw00244;
  wire nw00245;
  wire nw00246;
  wire nw00247;
  wire nw00248;
  wire nw00249;
  wire nw00250;
  wire nw00251;
  wire nw00252;
  wire nw00253;
  wire nw00254;
  wire nw00255;
  wire nw00256;
  wire nw00257;
  wire nw00258;
  wire nw00259;
  wire nw00260;
  wire nw00261;
  wire nw00262;
  wire nw00263;
  wire nw00264;
  wire nw00265;
  wire nw00266;
  wire nw00267;
  wire nw00268;
  wire nw00269;
  wire nw00270;
  wire nw00271;
  wire nw00272;
  wire nw00273;
  wire nw00274;
  wire nw00275;
  wire nw00276;
  wire nw00277;
  wire nw00278;
  wire nw00279;
  wire nw00280;
  wire nw00281;
  wire nw00282;
  wire nw00283;
  wire nw00284;
  wire nw00285;
  wire nw00286;
  wire nw00287;
  wire nw00288;
  wire nw00289;
  wire nw00290;
  wire nw00291;
  wire nw00292;
  wire nw00293;
  wire nw00294;
  wire nw00295;
  wire nw00296;
  wire nw00297;
  wire nw00298;
  wire nw00299;
  wire nw00300;
  wire nw00301;
  wire nw00302;
  wire nw00303;
  wire nw00304;
  wire nw00305;
  wire nw00306;
  wire nw00307;
  wire nw00308;
  wire nw00309;
  wire nw00310;
  wire nw00311;
  wire nw00312;
  wire nw00313;
  wire nw00314;
  wire nw00315;
  wire nw00316;
  wire nw00317;
  wire nw00318;
  wire nw00319;
  wire nw00320;
  wire nw00321;
  wire nw00322;
  wire nw00323;
  wire nw00324;
  wire nw00325;
  wire nw00326;
  wire nw00327;
  wire nw00328;
  wire nw00329;
  wire nw00330;
  wire nw00331;
  wire nw00332;
  wire nw00333;
  wire nw00334;
  wire nw00335;
  wire nw00336;
  wire nw00337;
  wire nw00338;
  wire nw00339;
  wire nw00340;
  wire nw00341;
  wire nw00342;
  wire nw00343;
  wire nw00344;
  wire nw00345;
  wire nw00346;
  wire nw00347;
  wire nw00348;
  wire nw00349;
  wire nw00350;
  wire nw00351;
  wire nw00352;
  wire nw00353;
  wire nw00354;
  wire nw00355;
  wire nw00356;
  wire nw00357;
  wire nw00358;
  wire nw00359;
  wire nw00360;
  wire nw00361;
  wire nw00362;
  wire nw00363;
  wire nw00364;
  wire nw00365;
  wire nw00366;
  wire nw00367;
  wire nw00368;
  wire nw00369;
  wire nw00370;
  wire nw00371;
  wire nw00372;
  wire nw00373;
  wire nw00374;
  wire nw00375;
  wire nw00376;
  wire nw00377;
  wire nw00378;
  wire nw00379;
  wire nw00380;
  wire nw00381;
  wire nw00382;
  wire nw00383;
  wire nw00384;
  wire nw00385;
  wire nw00386;
  wire nw00387;
  wire nw00388;
  wire nw00389;
  wire nw00390;
  wire nw00391;
  wire nw00392;
  wire nw00393;
  wire nw00394;
  wire nw00395;
  wire nw00396;
  wire nw00397;
  wire nw00398;
  wire nw00399;
  wire nw00400;
  wire nw00401;
  wire nw00402;
  wire nw00403;
  wire nw00404;
  wire nw00405;
  wire nw00406;
  wire nw00407;
  wire nw00408;
  wire nw00409;
  wire nw00410;
  wire nw00411;
  wire nw00412;
  wire nw00413;
  wire nw00414;
  wire nw00415;
  wire nw00416;
  wire nw00417;
  wire nw00418;
  wire nw00419;
  wire nw00420;
  wire nw00421;
  wire nw00422;
  wire nw00423;
  wire nw00424;
  wire nw00425;
  wire nw00426;
  wire nw00427;
  wire nw00428;
  wire nw00429;
  wire nw00430;
  wire nw00431;
  wire nw00432;
  wire nw00433;
  wire nw00434;
  wire nw00435;
  wire nw00436;
  wire nw00437;
  wire nw00438;
  wire nw00439;
  wire nw00440;
  wire nw00441;
  wire nw00442;
  wire nw00443;
  wire nw00444;
  wire nw00445;
  wire nw00446;
  wire nw00447;
  wire nw00448;
  wire nw00449;
  wire nw00450;
  wire nw00451;
  wire nw00452;
  wire nw00453;
  wire nw00454;
  wire nw00455;
  wire nw00456;
  wire nw00457;
  wire nw00458;
  wire nw00459;
  wire nw00460;
  wire nw00461;
  wire nw00462;
  wire nw00463;
  wire nw00464;
  wire nw00465;
  wire nw00466;
  wire nw00467;
  wire nw00468;
  wire nw00469;
  wire nw00470;
  wire nw00471;
  wire nw00472;
  wire nw00473;
  wire nw00474;
  wire nw00475;
  wire nw00476;
  wire nw00477;
  wire nw00478;
  wire nw00479;
  wire nw00480;
  wire nw00481;
  wire nw00482;
  wire nw00483;
  wire nw00484;
  wire nw00485;
  wire nw00486;
  wire nw00487;
  wire nw00488;
  wire nw00489;
  wire nw00490;
  wire nw00491;
  wire nw00492;
  wire nw00493;
  wire nw00494;
  wire nw00495;
  wire nw00496;
  wire nw00497;
  wire nw00498;
  wire nw00499;
  wire nw00500;
  wire nw00501;
  wire nw00502;
  wire nw00503;
  wire nw00504;
  wire nw00505;
  wire nw00506;
  wire nw00507;
  wire nw00508;
  wire nw00509;
  wire nw00510;
  wire nw00511;
  wire nw00512;
  wire nw00513;
  wire nw00514;
  wire nw00515;
  wire nw00516;
  wire nw00517;
  wire nw00518;
  wire nw00519;
  wire nw00520;
  wire nw00521;
  wire nw00522;
  wire nw00523;
  wire nw00524;
  wire nw00525;
  wire nw00526;
  wire nw00527;
  wire nw00528;
  wire nw00529;
  wire nw00530;
  wire nw00531;
  wire nw00532;
  wire nw00533;
  wire nw00534;
  wire nw00535;
  wire nw00536;
  wire nw00537;
  wire nw00538;
  wire nw00539;
  wire nw00540;
  wire nw00541;
  wire nw00542;
  wire nw00543;
  wire nw00544;
  wire nw00545;
  wire nw00546;
  wire nw00547;
  wire nw00548;
  wire nw00549;
  wire nw00550;
  wire nw00551;
  wire nw00552;
  wire nw00553;
  wire nw00554;
  wire nw00555;
  wire nw00556;
  wire nw00557;
  wire nw00558;
  wire nw00559;
  wire nw00560;
  wire nw00561;
  wire nw00562;
  wire nw00563;
  wire nw00564;
  wire nw00565;
  wire nw00566;
  wire nw00567;
  wire nw00568;
  wire nw00569;
  wire nw00570;
  wire nw00571;
  wire nw00572;
  wire nw00573;
  wire nw00574;
  wire nw00575;
  wire nw00576;
  wire nw00577;
  wire nw00578;
  wire nw00579;
  wire nw00580;
  wire nw00581;
  wire nw00582;
  wire nw00583;
  wire nw00584;
  wire nw00585;
  wire nw00586;
  wire nw00587;
  wire nw00588;
  wire nw00589;
  wire nw00590;
  wire nw00591;
  wire nw00592;
  wire nw00593;
  wire nw00594;
  wire nw00595;
  wire nw00596;
  wire nw00597;
  wire nw00598;
  wire nw00599;
  wire nw00600;
  wire nw00601;
  wire nw00602;
  wire nw00603;
  wire nw00604;
  wire nw00605;
  wire nw00606;
  wire nw00607;
  wire nw00608;
  wire nw00609;
  wire nw00610;
  wire nw00611;
  wire nw00612;
  wire nw00613;
  wire nw00614;
  wire nw00615;
  wire nw00616;
  wire nw00617;
  wire nw00618;
  wire nw00619;
  wire nw00620;
  wire nw00621;
  wire nw00622;
  wire nw00623;
  wire nw00624;
  wire nw00625;
  wire nw00626;
  wire nw00627;
  wire nw00628;
  wire nw00629;
  wire nw00630;
  wire nw00631;
  wire nw00632;
  wire nw00633;
  wire nw00634;
  wire nw00635;
  wire nw00636;
  wire nw00637;
  wire nw00638;
  wire nw00639;
  wire nw00640;
  wire nw00641;
  wire nw00642;
  wire nw00643;
  wire nw00644;
  wire nw00645;
  wire nw00646;
  wire nw00647;
  wire nw00648;
  wire nw00649;
  wire nw00650;
  wire nw00651;
  wire nw00652;
  wire nw00653;
  wire nw00654;
  wire nw00655;
  wire nw00656;
  wire nw00657;
  wire nw00658;
  wire nw00659;
  wire nw00660;
  wire nw00661;
  wire nw00662;
  wire nw00663;
  wire nw00664;
  wire nw00665;
  wire nw00666;
  wire nw00667;
  wire nw00668;
  wire nw00669;
  wire nw00670;
  wire nw00671;
  wire nw00672;
  wire nw00673;
  wire nw00674;
  wire nw00675;
  wire nw00676;
  wire nw00677;
  wire nw00678;
  wire nw00679;
  wire nw00680;
  wire nw00681;
  wire nw00682;
  wire nw00683;
  wire nw00684;
  wire nw00685;
  wire nw00686;
  wire nw00687;
  wire nw00688;
  wire nw00689;
  wire nw00690;
  wire nw00691;
  wire nw00692;
  wire nw00693;
  wire nw00694;
  wire nw00695;
  wire nw00696;
  wire nw00697;
  wire nw00698;
  wire nw00699;
  wire nw00700;
  wire nw00701;
  wire nw00702;
  wire nw00703;
  wire nw00704;
  wire nw00705;
  wire nw00706;
  wire nw00707;
  wire nw00708;
  wire nw00709;
  wire nw00710;
  wire nw00711;
  wire nw00712;
  wire nw00713;
  wire nw00714;
  wire nw00715;
  wire nw00716;
  wire nw00717;
  wire nw00718;
  wire nw00719;
  wire nw00720;
  wire nw00721;
  wire nw00722;
  wire nw00723;
  wire nw00724;
  wire nw00725;
  wire nw00726;
  wire nw00727;
  wire nw00728;
  wire nw00729;
  wire nw00730;
  wire nw00731;
  wire nw00732;
  wire nw00733;
  wire nw00734;
  wire nw00735;
  wire nw00736;
  wire nw00737;
  wire nw00738;
  wire nw00739;
  wire nw00740;
  wire nw00741;
  wire nw00742;
  wire nw00743;
  wire nw00744;
  wire nw00745;
  wire nw00746;
  wire nw00747;
  wire nw00748;
  wire nw00749;
  wire nw00750;
  wire nw00751;
  wire nw00752;
  wire nw00753;
  wire nw00754;
  wire nw00755;
  wire nw00756;
  wire nw00757;
  wire nw00758;
  wire nw00759;
  wire nw00760;
  wire nw00761;
  wire nw00762;
  wire nw00763;
  wire nw00764;
  wire nw00765;
  wire nw00766;
  wire nw00767;
  wire nw00768;
  wire nw00769;
  wire nw00770;
  wire nw00771;
  wire nw00772;
  wire nw00773;
  wire nw00774;
  wire nw00775;
  wire nw00776;
  wire nw00777;
  wire nw00778;
  wire nw00779;
  wire nw00780;
  wire nw00781;
  wire nw00782;
  wire nw00783;
  wire nw00784;
  wire nw00785;
  wire nw00786;
  wire nw00787;
  wire nw00788;
  wire nw00789;
  wire nw00790;
  wire nw00791;
  wire nw00792;
  wire nw00793;
  wire nw00794;
  wire nw00795;
  wire nw00796;
  wire nw00797;
  wire nw00798;
  wire nw00799;
  wire nw00800;
  wire nw00801;
  wire nw00802;
  wire nw00803;
  wire nw00804;
  wire nw00805;
  wire nw00806;
  wire nw00807;
  wire nw00808;
  wire nw00809;
  wire nw00810;
  wire nw00811;
  wire nw00812;
  wire nw00813;
  wire nw00814;
  wire nw00815;
  wire nw00816;
  wire nw00817;
  wire nw00818;
  wire nw00819;
  wire nw00820;
  wire nw00821;
  wire nw00822;
  wire nw00823;
  wire nw00824;
  wire nw00825;
  wire nw00826;
  wire nw00827;
  wire nw00828;
  wire nw00829;
  wire nw00830;
  wire nw00831;
  wire nw00832;
  wire nw00833;
  wire nw00834;
  wire nw00835;
  wire nw00836;
  wire nw00837;
  wire nw00838;
  wire nw00839;
  wire nw00840;
  wire nw00841;
  wire nw00842;
  wire nw00843;
  wire nw00844;
  wire nw00845;
  wire nw00846;
  wire nw00847;
  wire nw00848;
  wire nw00849;
  wire nw00850;
  wire nw00851;
  wire nw00852;
  wire nw00853;
  wire nw00854;
  wire nw00855;
  wire nw00856;
  wire nw00857;
  wire nw00858;
  wire nw00859;
  wire nw00860;
  wire nw00861;
  wire nw00862;
  wire nw00863;
  wire nw00864;
  wire nw00865;
  wire nw00866;
  wire nw00867;
  wire nw00868;
  wire nw00869;
  wire nw00870;
  wire nw00871;
  wire nw00872;
  wire nw00873;
  wire nw00874;
  wire nw00875;
  wire nw00876;
  wire nw00877;
  wire nw00878;
  wire nw00879;
  wire nw00880;
  wire nw00881;
  wire nw00882;
  wire nw00883;
  wire nw00884;
  wire nw00885;
  wire nw00886;
  wire nw00887;
  wire nw00888;
  wire nw00889;
  wire nw00890;
  wire nw00891;
  wire nw00892;
  wire nw00893;
  wire nw00894;
  wire nw00895;
  wire nw00896;
  wire nw00897;
  wire nw00898;
  wire nw00899;
  wire nw00900;
  wire nw00901;
  wire nw00902;
  wire nw00903;
  wire nw00904;
  wire nw00905;
  wire nw00906;
  wire nw00907;
  wire nw00908;
  wire nw00909;
  wire nw00910;
  wire nw00911;
  wire nw00912;
  wire nw00913;
  wire nw00914;
  wire nw00915;
  wire nw00916;
  wire nw00917;
  wire nw00918;
  wire nw00919;
  wire nw00920;
  wire nw00921;
  wire nw00922;
  wire nw00923;
  wire nw00924;
  wire nw00925;
  wire nw00926;
  wire nw00927;
  wire nw00928;
  wire nw00929;
  wire nw00930;
  wire nw00931;
  wire nw00932;
  wire nw00933;
  wire nw00934;
  wire nw00935;
  wire nw00936;
  wire nw00937;
  wire nw00938;
  wire nw00939;
  wire nw00940;
  wire nw00941;
  wire nw00942;
  wire nw00943;
  wire nw00944;
  wire nw00945;
  wire nw00946;
  wire nw00947;
  wire nw00948;
  wire nw00949;
  wire nw00950;
  wire nw00951;
  wire nw00952;
  wire nw00953;
  wire nw00954;
  wire nw00955;
  wire nw00956;
  wire nw00957;
  wire nw00958;
  wire nw00959;
  wire nw00960;
  wire nw00961;
  wire nw00962;
  wire nw00963;
  wire nw00964;
  wire nw00965;
  wire nw00966;
  wire nw00967;
  wire nw00968;
  wire nw00969;
  wire nw00970;
  wire nw00971;
  wire nw00972;
  wire nw00973;
  wire nw00974;
  wire nw00975;
  wire nw00976;
  wire nw00977;
  wire nw00978;
  wire nw00979;
  wire nw00980;
  wire nw00981;
  wire nw00982;
  wire nw00983;
  wire nw00984;
  wire nw00985;
  wire nw00986;
  wire nw00987;
  wire nw00988;
  wire nw00989;
  wire nw00990;
  wire nw00991;
  wire nw00992;
  wire nw00993;
  wire nw00994;
  wire nw00995;
  wire nw00996;
  wire nw00997;
  wire nw00998;
  wire nw00999;
  wire nw01000;
  wire nw01001;
  wire nw01002;
  wire nw01003;
  wire nw01004;
  wire nw01005;
  wire nw01006;
  wire nw01007;
  wire nw01008;
  wire nw01009;
  wire nw01010;
  wire nw01011;
  wire nw01012;
  wire nw01013;
  wire nw01014;
  wire nw01015;
  wire nw01016;
  wire nw01017;
  wire nw01018;
  wire nw01019;
  wire nw01020;
  wire nw01021;
  wire nw01022;
  wire nw01023;
  wire nw01024;
  wire nw01025;
  wire nw01026;
  wire nw01027;
  wire nw01028;
  wire nw01029;
  wire nw01030;
  wire nw01031;
  wire nw01032;
  wire nw01033;
  wire nw01034;
  wire nw01035;
  wire nw01036;
  wire nw01037;
  wire nw01038;
  wire nw01039;
  wire nw01040;
  wire nw01041;
  wire nw01042;
  wire nw01043;
  wire nw01044;
  wire nw01045;
  wire nw01046;
  wire nw01047;
  wire nw01048;
  wire nw01049;
  wire nw01050;
  wire nw01051;
  wire nw01052;
  wire nw01053;
  wire nw01054;
  wire nw01055;
  wire nw01056;
  wire nw01057;
  wire nw01058;
  wire nw01059;
  wire nw01060;
  wire nw01061;
  wire nw01062;
  wire nw01063;
  wire nw01064;
  wire nw01065;
  wire nw01066;
  wire nw01067;
  wire nw01068;
  wire nw01069;
  wire nw01070;
  wire nw01071;
  wire nw01072;
  wire nw01073;
  wire nw01074;
  wire nw01075;
  wire nw01076;
  wire nw01077;
  wire nw01078;
  wire nw01079;
  wire nw01080;
  wire nw01081;
  wire nw01082;
  wire nw01083;
  wire nw01084;
  wire nw01085;
  wire nw01086;
  wire nw01087;
  wire nw01088;
  wire nw01089;
  wire nw01090;
  wire nw01091;
  wire nw01092;
  wire nw01093;
  wire nw01094;
  wire nw01095;
  wire nw01096;
  wire nw01097;
  wire nw01098;
  wire nw01099;
  wire nw01100;
  wire nw01101;
  wire nw01102;
  wire nw01103;
  wire nw01104;
  wire nw01105;
  wire nw01106;
  wire nw01107;
  wire nw01108;
  wire nw01109;
  wire nw01110;
  wire nw01111;
  wire nw01112;
  wire nw01113;
  wire nw01114;
  wire nw01115;
  wire nw01116;
  wire nw01117;
  wire nw01118;
  wire nw01119;
  wire nw01120;
  wire nw01121;
  wire nw01122;
  wire nw01123;
  wire nw01124;
  wire nw01125;
  wire nw01126;
  wire nw01127;
  wire nw01128;
  wire nw01129;
  wire nw01130;
  wire nw01131;
  wire nw01132;
  wire nw01133;
  wire nw01134;
  wire nw01135;
  wire nw01136;
  wire nw01137;
  wire nw01138;
  wire nw01139;
  wire nw01140;
  wire nw01141;
  wire nw01142;
  wire nw01143;
  wire nw01144;
  wire nw01145;
  wire nw01146;
  wire nw01147;
  wire nw01148;
  wire nw01149;
  wire nw01150;
  wire nw01151;
  wire nw01152;
  wire nw01153;
  wire nw01154;
  wire nw01155;
  wire nw01156;
  wire nw01157;
  wire nw01158;
  wire nw01159;
  wire nw01160;
  wire nw01161;
  wire nw01162;
  wire nw01163;
  wire nw01164;
  wire nw01165;
  wire nw01166;
  wire nw01167;
  wire nw01168;
  wire nw01169;
  wire nw01170;
  wire nw01171;
  wire nw01172;
  wire nw01173;
  wire nw01174;
  wire nw01175;
  wire nw01176;
  wire nw01177;
  wire nw01178;
  wire nw01179;
  wire nw01180;
  wire nw01181;
  wire nw01182;
  wire nw01183;
  wire nw01184;
  wire nw01185;
  wire nw01186;
  wire nw01187;
  wire nw01188;
  wire nw01189;
  wire nw01190;
  wire nw01191;
  wire nw01192;
  wire nw01193;
  wire nw01194;
  wire nw01195;
  wire nw01196;
  wire nw01197;
  wire nw01198;
  wire nw01199;
  wire nw01200;
  wire nw01201;
  wire nw01202;
  wire nw01203;
  wire nw01204;
  wire nw01205;
  wire nw01206;
  wire nw01207;
  wire nw01208;
  wire nw01209;
  wire nw01210;
  wire nw01211;
  wire nw01212;
  wire nw01213;
  wire nw01214;
  wire nw01215;
  wire nw01216;
  wire nw01217;
  wire nw01218;
  wire nw01219;
  wire nw01220;
  wire nw01221;
  wire nw01222;
  wire nw01223;
  wire nw01224;
  wire nw01225;
  wire nw01226;
  wire nw01227;
  wire nw01228;
  wire nw01229;
  wire nw01230;
  wire nw01231;
  wire nw01232;
  wire nw01233;
  wire nw01234;
  wire nw01235;
  wire nw01236;
  wire nw01237;
  wire nw01238;
  wire nw01239;
  wire nw01240;
  wire nw01241;
  wire nw01242;
  wire nw01243;
  wire nw01244;
  wire nw01245;
  wire nw01246;
  wire nw01247;
  wire nw01248;
  wire nw01249;
  wire nw01250;
  wire nw01251;
  wire nw01252;
  wire nw01253;
  wire nw01254;
  wire nw01255;
  wire nw01256;
  wire nw01257;
  wire nw01258;
  wire nw01259;
  wire nw01260;
  wire nw01261;
  wire nw01262;
  wire nw01263;
  wire nw01264;
  wire nw01265;
  wire nw01266;
  wire nw01267;
  wire nw01268;
  wire nw01269;
  wire nw01270;
  wire nw01271;
  wire nw01272;
  wire nw01273;
  wire nw01274;
  wire nw01275;
  wire nw01276;
  wire nw01277;
  wire nw01278;
  wire nw01279;
  wire nw01280;
  wire nw01281;
  wire nw01282;
  wire nw01283;
  wire nw01284;
  wire nw01285;
  wire nw01286;
  wire nw01287;
  wire nw01288;
  wire nw01289;
  wire nw01290;
  wire nw01291;
  wire nw01292;
  wire nw01293;
  wire nw01294;
  wire nw01295;
  wire nw01296;
  wire nw01297;
  wire nw01298;
  wire nw01299;
  wire nw01300;
  wire nw01301;
  wire nw01302;
  wire nw01303;
  wire nw01304;
  wire nw01305;
  wire nw01306;
  wire nw01307;
  wire nw01308;
  wire nw01309;
  wire nw01310;
  wire nw01311;
  wire nw01312;
  wire nw01313;
  wire nw01314;
  wire nw01315;
  wire nw01316;
  wire nw01317;
  wire nw01318;
  wire nw01319;
  wire nw01320;
  wire nw01321;
  wire nw01322;
  wire nw01323;
  wire nw01324;
  wire nw01325;
  wire nw01326;
  wire nw01327;
  wire nw01328;
  wire nw01329;
  wire nw01330;
  wire nw01331;
  wire nw01332;
  wire nw01333;
  wire nw01334;
  wire nw01335;
  wire nw01336;
  wire nw01337;
  wire nw01338;
  wire nw01339;
  wire nw01340;
  wire nw01341;
  wire nw01342;
  wire nw01343;
  wire nw01344;
  wire nw01345;
  wire nw01346;
  wire nw01347;
  wire nw01348;
  wire nw01349;
  wire nw01350;
  wire nw01351;
  wire nw01352;
  wire nw01353;
  wire nw01354;
  wire nw01355;
  wire nw01356;
  wire nw01357;
  wire nw01358;
  wire nw01359;
  wire nw01360;
  wire nw01361;
  wire nw01362;
  wire nw01363;
  wire nw01364;
  wire nw01365;
  wire nw01366;
  wire nw01367;
  wire nw01368;
  wire nw01369;
  wire nw01370;
  wire nw01371;
  wire nw01372;
  wire nw01373;
  wire nw01374;
  wire nw01375;
  wire nw01376;
  wire nw01377;
  wire nw01378;
  wire nw01379;
  wire nw01380;
  wire nw01381;
  wire nw01382;
  wire nw01383;
  wire nw01384;
  wire nw01385;
  wire nw01386;
  wire nw01387;
  wire nw01388;
  wire nw01389;
  wire nw01390;
  wire nw01391;
  wire nw01392;
  wire nw01393;
  wire nw01394;
  wire nw01395;
  wire nw01396;
  wire nw01397;
  wire nw01398;
  wire nw01399;
  wire nw01400;
  wire nw01401;
  wire nw01402;
  wire nw01403;
  wire nw01404;
  wire nw01405;
  wire nw01406;
  wire nw01407;
  wire nw01408;
  wire nw01409;
  wire nw01410;
  wire nw01411;
  wire nw01412;
  wire nw01413;
  wire nw01414;
  wire nw01415;
  wire nw01416;
  wire nw01417;
  wire nw01418;
  wire nw01419;
  wire nw01420;
  wire nw01421;
  wire nw01422;
  wire nw01423;
  wire nw01424;
  wire nw01425;
  wire nw01426;
  wire nw01427;
  wire nw01428;
  wire nw01429;
  wire nw01430;
  wire nw01431;
  wire nw01432;
  wire nw01433;
  wire nw01434;
  wire nw01435;
  wire nw01436;
  wire nw01437;
  wire nw01438;
  wire nw01439;
  wire nw01440;
  wire nw01441;
  wire nw01442;
  wire nw01443;
  wire nw01444;
  wire nw01445;
  wire nw01446;
  wire nw01447;
  wire nw01448;
  wire nw01449;
  wire nw01450;
  wire nw01451;
  wire nw01452;
  wire nw01453;
  wire nw01454;
  wire nw01455;
  wire nw01456;
  wire nw01457;
  wire nw01458;
  wire nw01459;
  wire nw01460;
  wire nw01461;
  wire nw01462;
  wire nw01463;
  wire nw01464;
  wire nw01465;
  wire nw01466;
  wire nw01467;
  wire nw01468;
  wire nw01469;
  wire nw01470;
  wire nw01471;
  wire nw01472;
  wire nw01473;
  wire nw01474;
  wire nw01475;
  wire nw01476;
  wire nw01477;
  wire nw01478;
  wire nw01479;
  wire nw01480;
  wire nw01481;
  wire nw01482;
  wire nw01483;
  wire nw01484;
  wire nw01485;
  wire nw01486;
  wire nw01487;
  wire nw01488;
  wire nw01489;
  wire nw01490;
  wire nw01491;
  wire nw01492;
  wire nw01493;
  wire nw01494;
  wire nw01495;
  wire nw01496;
  wire nw01497;
  wire nw01498;
  wire nw01499;
  wire nw01500;
  wire nw01501;
  wire nw01502;
  wire nw01503;
  wire nw01504;
  wire nw01505;
  wire nw01506;
  wire nw01507;
  wire nw01508;
  wire nw01509;
  wire nw01510;
  wire nw01511;
  wire nw01512;
  wire nw01513;
  wire nw01514;
  wire nw01515;
  wire nw01516;
  wire nw01517;
  wire nw01518;
  wire nw01519;
  wire nw01520;
  wire nw01521;
  wire nw01522;
  wire nw01523;
  wire nw01524;
  wire nw01525;
  wire nw01526;
  wire nw01527;
  wire nw01528;
  wire nw01529;
  wire nw01530;
  wire nw01531;
  wire nw01532;
  wire nw01533;
  wire nw01534;
  wire nw01535;
  wire nw01536;
  wire nw01537;
  wire nw01538;
  wire nw01539;
  wire nw01540;
  wire nw01541;
  wire nw01542;
  wire nw01543;
  wire nw01544;
  wire nw01545;
  wire nw01546;
  wire nw01547;
  wire nw01548;
  wire nw01549;
  wire nw01550;
  wire nw01551;
  wire nw01552;
  wire nw01553;
  wire nw01554;
  wire nw01555;
  wire nw01556;
  wire nw01557;
  wire nw01558;
  wire nw01559;
  wire nw01560;
  wire nw01561;
  wire nw01562;
  wire nw01563;
  wire nw01564;
  wire nw01565;
  wire nw01566;
  wire nw01567;
  wire nw01568;
  wire nw01569;
  wire nw01570;
  wire nw01571;
  wire nw01572;
  wire nw01573;
  wire nw01574;
  wire nw01575;
  wire nw01576;
  wire nw01577;
  wire nw01578;
  wire nw01579;
  wire nw01580;
  wire nw01581;
  wire nw01582;
  wire nw01583;
  wire nw01584;
  wire nw01585;
  wire nw01586;
  wire nw01587;
  wire nw01588;
  wire nw01589;
  wire nw01590;
  wire nw01591;
  wire nw01592;
  wire nw01593;
  wire nw01594;
  wire nw01595;
  wire nw01596;
  wire nw01597;
  wire nw01598;
  wire nw01599;
  wire nw01600;
  wire nw01601;
  wire nw01602;
  wire nw01603;
  wire nw01604;
  wire nw01605;
  wire nw01606;
  wire nw01607;
  wire nw01608;
  wire nw01609;
  wire nw01610;
  wire nw01611;
  wire nw01612;
  wire nw01613;
  wire nw01614;
  wire nw01615;
  wire nw01616;
  wire nw01617;
  wire nw01618;
  wire nw01619;
  wire nw01620;
  wire nw01621;
  wire nw01622;
  wire nw01623;
  wire nw01624;
  wire nw01625;
  wire nw01626;
  wire nw01627;
  wire nw01628;
  wire nw01629;
  wire nw01630;
  wire nw01631;
  wire nw01632;
  wire nw01633;
  wire nw01634;
  wire nw01635;
  wire nw01636;
  wire nw01637;
  wire nw01638;
  wire nw01639;
  wire nw01640;
  wire nw01641;
  wire nw01642;
  wire nw01643;
  wire nw01644;
  wire nw01645;
  wire nw01646;
  wire nw01647;
  wire nw01648;
  wire nw01649;
  wire nw01650;
  wire nw01651;
  wire nw01652;
  wire nw01653;
  wire nw01654;
  wire nw01655;
  wire nw01656;
  wire nw01657;
  wire nw01658;
  wire nw01659;
  wire nw01660;
  wire nw01661;
  wire nw01662;
  wire nw01663;
  wire nw01664;
  wire nw01665;
  wire nw01666;
  wire nw01667;
  wire nw01668;
  wire nw01669;
  wire nw01670;
  wire nw01671;
  wire nw01672;
  wire nw01673;
  wire nw01674;
  wire nw01675;
  wire nw01676;
  wire nw01677;
  wire nw01678;
  wire nw01679;
  wire nw01680;
  wire nw01681;
  wire nw01682;
  wire nw01683;
  wire nw01684;
  wire nw01685;
  wire nw01686;
  wire nw01687;
  wire nw01688;
  wire nw01689;
  wire nw01690;
  wire nw01691;
  wire nw01692;
  wire nw01693;
  wire nw01694;
  wire nw01695;
  wire nw01696;
  wire nw01697;
  wire nw01698;
  wire nw01699;
  wire nw01700;
  wire nw01701;
  wire nw01702;
  wire nw01703;
  wire nw01704;
  wire nw01705;
  wire nw01706;
  wire nw01707;
  wire nw01708;
  wire nw01709;
  wire nw01710;
  wire nw01711;
  wire nw01712;
  wire nw01713;
  wire nw01714;
  wire nw01715;
  wire nw01716;
  wire nw01717;
  wire nw01718;
  wire nw01719;
  wire nw01720;
  wire nw01721;
  wire nw01722;
  wire nw01723;
  wire nw01724;
  wire nw01725;
  wire nw01726;
  wire nw01727;
  wire nw01728;
  wire nw01729;
  wire nw01730;
  wire nw01731;
  wire nw01732;
  wire nw01733;
  wire nw01734;
  wire nw01735;
  wire nw01736;
  wire nw01737;
  wire nw01738;
  wire nw01739;
  wire nw01740;
  wire nw01741;
  wire nw01742;
  wire nw01743;
  wire nw01744;
  wire nw01745;
  wire nw01746;
  wire nw01747;
  wire nw01748;
  wire nw01749;
  wire nw01750;
  wire nw01751;
  wire nw01752;
  wire nw01753;
  wire nw01754;
  wire nw01755;
  wire nw01756;
  wire nw01757;
  wire nw01758;
  wire nw01759;
  wire nw01760;
  wire nw01761;
  wire nw01762;
  wire nw01763;
  wire nw01764;
  wire nw01765;
  wire nw01766;
  wire nw01767;
  wire nw01768;
  wire nw01769;
  wire nw01770;
  wire nw01771;
  wire nw01772;
  wire nw01773;
  wire nw01774;
  wire nw01775;
  wire nw01776;
  wire nw01777;
  wire nw01778;
  wire nw01779;
  wire nw01780;
  wire nw01781;
  wire nw01782;
  wire nw01783;
  wire nw01784;
  wire nw01785;
  wire nw01786;
  wire nw01787;
  wire nw01788;
  wire nw01789;
  wire nw01790;
  wire nw01791;
  wire nw01792;
  wire nw01793;
  wire nw01794;
  wire nw01795;
  wire nw01796;
  wire nw01797;
  wire nw01798;
  wire nw01799;
  wire nw01800;
  wire nw01801;
  wire nw01802;
  wire nw01803;
  wire nw01804;
  wire nw01805;
  wire nw01806;
  wire nw01807;
  wire nw01808;
  wire nw01809;
  wire nw01810;
  wire nw01811;
  wire nw01812;
  wire nw01813;
  wire nw01814;
  wire nw01815;
  wire nw01816;
  wire nw01817;
  wire nw01818;
  wire nw01819;
  wire nw01820;
  wire nw01821;
  wire nw01822;
  wire nw01823;
  wire nw01824;
  wire nw01825;
  wire nw01826;
  wire nw01827;
  wire nw01828;
  wire nw01829;
  wire nw01830;
  wire nw01831;
  wire nw01832;
  wire nw01833;
  wire nw01834;
  wire nw01835;
  wire nw01836;
  wire nw01837;
  wire nw01838;
  wire nw01839;
  wire nw01840;
  wire nw01841;
  wire nw01842;
  wire nw01843;
  wire nw01844;
  wire nw01845;
  wire nw01846;
  wire nw01847;
  wire nw01848;
  wire nw01849;
  wire nw01850;
  wire nw01851;
  wire nw01852;
  wire nw01853;
  wire nw01854;
  wire nw01855;
  wire nw01856;
  wire nw01857;
  wire nw01858;
  wire nw01859;
  wire nw01860;
  wire nw01861;
  wire nw01862;
  wire nw01863;
  wire nw01864;
  wire nw01865;
  wire nw01866;
  wire nw01867;
  wire nw01868;
  wire nw01869;
  wire nw01870;
  wire nw01871;
  wire nw01872;
  wire nw01873;
  wire nw01874;
  wire nw01875;
  wire nw01876;
  wire nw01877;
  wire nw01878;
  wire nw01879;
  wire nw01880;
  wire nw01881;
  wire nw01882;
  wire nw01883;
  wire nw01884;
  wire nw01885;
  wire nw01886;
  wire nw01887;
  wire nw01888;
  wire nw01889;
  wire nw01890;
  wire nw01891;
  wire nw01892;
  wire nw01893;
  wire nw01894;
  wire nw01895;
  wire nw01896;
  wire nw01897;
  wire nw01898;
  wire nw01899;
  wire nw01900;
  wire nw01901;
  wire nw01902;
  wire nw01903;
  wire nw01904;
  wire nw01905;
  wire nw01906;
  wire nw01907;
  wire nw01908;
  wire nw01909;
  wire nw01910;
  wire nw01911;
  wire nw01912;
  wire nw01913;
  wire nw01914;
  wire nw01915;
  wire nw01916;
  wire nw01917;
  wire nw01918;
  wire nw01919;
  wire nw01920;
  wire nw01921;
  wire nw01922;
  wire nw01923;
  wire nw01924;
  wire nw01925;
  wire nw01926;
  wire nw01927;
  wire nw01928;
  wire nw01929;
  wire nw01930;
  wire nw01931;
  wire nw01932;
  wire nw01933;
  wire nw01934;
  wire nw01935;
  wire nw01936;
  wire nw01937;
  wire nw01938;
  wire nw01939;
  wire nw01940;
  wire nw01941;
  wire nw01942;
  wire nw01943;
  wire nw01944;
  wire nw01945;
  wire nw01946;
  wire nw01947;
  wire nw01948;
  wire nw01949;
  wire nw01950;
  wire nw01951;
  wire nw01952;
  wire nw01953;
  wire nw01954;
  wire nw01955;
  wire nw01956;
  wire nw01957;
  wire nw01958;
  wire nw01959;
  wire nw01960;
  wire nw01961;
  wire nw01962;
  wire nw01963;
  wire nw01964;
  wire nw01965;
  wire nw01966;
  wire nw01967;
  wire nw01968;
  wire nw01969;
  wire nw01970;
  wire nw01971;
  wire nw01972;
  wire nw01973;
  wire nw01974;
  wire nw01975;
  wire nw01976;
  wire nw01977;
  wire nw01978;
  wire nw01979;
  wire nw01980;
  wire nw01981;
  wire nw01982;
  wire nw01983;
  wire nw01984;
  wire nw01985;
  wire nw01986;
  wire nw01987;
  wire nw01988;
  wire nw01989;
  wire nw01990;
  wire nw01991;
  wire nw01992;
  wire nw01993;
  wire nw01994;
  wire nw01995;
  wire nw01996;
  wire nw01997;
  wire nw01998;
  wire nw01999;
  wire nw02000;
  wire nw02001;
  wire nw02002;
  wire nw02003;
  wire nw02004;
  wire nw02005;
  wire nw02006;
  wire nw02007;
  wire nw02008;
  wire nw02009;
  wire nw02010;
  wire nw02011;
  wire nw02012;
  wire nw02013;
  wire nw02014;
  wire nw02015;
  wire nw02016;
  wire nw02017;
  wire nw02018;
  wire nw02019;
  wire nw02020;
  wire nw02021;
  wire nw02022;
  wire nw02023;
  wire nw02024;
  wire nw02025;
  wire nw02026;
  wire nw02027;
  wire nw02028;
  wire nw02029;
  wire nw02030;
  wire nw02031;
  wire nw02032;
  wire nw02033;
  wire nw02034;
  wire nw02035;
  wire nw02036;
  wire nw02037;
  wire nw02038;
  wire nw02039;
  wire nw02040;
  wire nw02041;
  wire nw02042;
  wire nw02043;
  wire nw02044;
  wire nw02045;
  wire nw02046;
  wire nw02047;
  wire nw02048;
  wire nw02049;
  wire nw02050;
  wire nw02051;
  wire nw02052;
  wire nw02053;
  wire nw02054;
  wire nw02055;
  wire nw02056;
  wire nw02057;
  wire nw02058;
  wire nw02059;
  wire nw02060;
  wire nw02061;
  wire nw02062;
  wire nw02063;
  wire nw02064;
  wire nw02065;
  wire nw02066;
  wire nw02067;
  wire nw02068;
  wire nw02069;
  wire nw02070;
  wire nw02071;
  wire nw02072;
  wire nw02073;
  wire nw02074;
  wire nw02075;
  wire nw02076;
  wire nw02077;
  wire nw02078;
  wire nw02079;
  wire nw02080;
  wire nw02081;
  wire nw02082;
  wire nw02083;
  wire nw02084;
  wire nw02085;
  wire nw02086;
  wire nw02087;
  wire nw02088;
  wire nw02089;
  wire nw02090;
  wire nw02091;
  wire nw02092;
  wire nw02093;
  wire nw02094;
  wire nw02095;
  wire nw02096;
  wire nw02097;
  wire nw02098;
  wire nw02099;
  wire nw02100;
  wire nw02101;
  wire nw02102;
  wire nw02103;
  wire nw02104;
  wire nw02105;
  wire nw02106;
  wire nw02107;
  wire nw02108;
  wire nw02109;
  wire nw02110;
  wire nw02111;
  wire nw02112;
  wire nw02113;
  wire nw02114;
  wire nw02115;
  wire nw02116;
  wire nw02117;
  wire nw02118;
  wire nw02119;
  wire nw02120;
  wire nw02121;
  wire nw02122;
  wire nw02123;
  wire nw02124;
  wire nw02125;
  wire nw02126;
  wire nw02127;
  wire nw02128;
  wire nw02129;
  wire nw02130;
  wire nw02131;
  wire nw02132;
  wire nw02133;
  wire nw02134;
  wire nw02135;
  wire nw02136;
  wire nw02137;
  wire nw02138;
  wire nw02139;
  wire nw02140;
  wire nw02141;
  wire nw02142;
  wire nw02143;
  wire nw02144;
  wire nw02145;
  wire nw02146;
  wire nw02147;
  wire nw02148;
  wire nw02149;
  wire nw02150;
  wire nw02151;
  wire nw02152;
  wire nw02153;
  wire nw02154;
  wire nw02155;
  wire nw02156;
  wire nw02157;
  wire nw02158;
  wire nw02159;
  wire nw02160;
  wire nw02161;
  wire nw02162;
  wire nw02163;
  wire nw02164;
  wire nw02165;
  wire nw02166;
  wire nw02167;
  wire nw02168;
  wire nw02169;
  wire nw02170;
  wire nw02171;
  wire nw02172;
  wire nw02173;
  wire nw02174;
  wire nw02175;
  wire nw02176;
  wire nw02177;
  wire nw02178;
  wire nw02179;
  wire nw02180;
  wire nw02181;
  wire nw02182;
  wire nw02183;
  wire nw02184;
  wire nw02185;
  wire nw02186;
  wire nw02187;
  wire nw02188;
  wire nw02189;
  wire nw02190;
  wire nw02191;
  wire nw02192;
  wire nw02193;
  wire nw02194;
  wire nw02195;
  wire nw02196;
  wire nw02197;
  wire nw02198;
  wire nw02199;
  wire nw02200;
  wire nw02201;
  wire nw02202;
  wire nw02203;
  wire nw02204;
  wire nw02205;
  wire nw02206;
  wire nw02207;
  wire nw02208;
  wire nw02209;
  wire nw02210;
  wire nw02211;
  wire nw02212;
  wire nw02213;
  wire nw02214;
  wire nw02215;
  wire nw02216;
  wire nw02217;
  wire nw02218;
  wire nw02219;
  wire nw02220;
  wire nw02221;
  wire nw02222;
  wire nw02223;
  wire nw02224;
  wire nw02225;
  wire nw02226;
  wire nw02227;
  wire nw02228;
  wire nw02229;
  wire nw02230;
  wire nw02231;
  wire nw02232;
  wire nw02233;
  wire nw02234;
  wire nw02235;
  wire nw02236;
  wire nw02237;
  wire nw02238;
  wire nw02239;
  wire nw02240;
  wire nw02241;
  wire nw02242;
  wire nw02243;
  wire nw02244;
  wire nw02245;
  wire nw02246;
  wire nw02247;
  wire nw02248;
  wire nw02249;
  wire nw02250;
  wire nw02251;
  wire nw02252;
  wire nw02253;
  wire nw02254;
  wire nw02255;
  wire nw02256;
  wire nw02257;
  wire nw02258;
  wire nw02259;
  wire nw02260;
  wire nw02261;
  wire nw02262;
  wire nw02263;
  wire nw02264;
  wire nw02265;
  wire nw02266;
  wire nw02267;
  wire nw02268;
  wire nw02269;
  wire nw02270;
  wire nw02271;
  wire nw02272;
  wire nw02273;
  wire nw02274;
  wire nw02275;
  wire nw02276;
  wire nw02277;
  wire nw02278;
  wire nw02279;
  wire nw02280;
  wire nw02281;
  wire nw02282;
  wire nw02283;
  wire nw02284;
  wire nw02285;
  wire nw02286;
  wire nw02287;
  wire nw02288;
  wire nw02289;
  wire nw02290;
  wire nw02291;
  wire nw02292;
  wire nw02293;
  wire nw02294;
  wire nw02295;
  wire nw02296;
  wire nw02297;
  wire nw02298;
  wire nw02299;
  wire nw02300;
  wire nw02301;
  wire nw02302;
  wire nw02303;
  wire nw02304;
  wire nw02305;
  wire nw02306;
  wire nw02307;
  wire nw02308;
  wire nw02309;
  wire nw02310;
  wire nw02311;
  wire nw02312;
  wire nw02313;
  wire nw02314;
  wire nw02315;
  wire nw02316;
  wire nw02317;
  wire nw02318;
  wire nw02319;
  wire nw02320;
  wire nw02321;
  wire nw02322;
  wire nw02323;
  wire nw02324;
  wire nw02325;
  wire nw02326;
  wire nw02327;
  wire nw02328;
  wire nw02329;
  wire nw02330;
  wire nw02331;
  wire nw02332;
  wire nw02333;
  wire nw02334;
  wire nw02335;
  wire nw02336;
  wire nw02337;
  wire nw02338;
  wire nw02339;
  wire nw02340;
  wire nw02341;
  wire nw02342;
  wire nw02343;
  wire nw02344;
  wire nw02345;
  wire nw02346;
  wire nw02347;
  wire nw02348;
  wire nw02349;
  wire nw02350;
  wire nw02351;
  wire nw02352;
  wire nw02353;
  wire nw02354;
  wire nw02355;
  wire nw02356;
  wire nw02357;
  wire nw02358;
  wire nw02359;
  wire nw02360;
  wire nw02361;
  wire nw02362;
  wire nw02363;
  wire nw02364;
  wire nw02365;
  wire nw02366;
  wire nw02367;
  wire nw02368;
  wire nw02369;
  wire nw02370;
  wire nw02371;
  wire nw02372;
  wire nw02373;
  wire nw02374;
  wire nw02375;
  wire nw02376;
  wire nw02377;
  wire nw02378;
  wire nw02379;
  wire nw02380;
  wire nw02381;
  wire nw02382;
  wire nw02383;
  wire nw02384;
  wire nw02385;
  wire nw02386;
  wire nw02387;
  wire nw02388;
  wire nw02389;
  wire nw02390;
  wire nw02391;
  wire nw02392;
  wire nw02393;
  wire nw02394;
  wire nw02395;
  wire nw02396;
  wire nw02397;
  wire nw02398;
  wire nw02399;
  wire nw02400;
  wire nw02401;
  wire nw02402;
  wire nw02403;
  wire nw02404;
  wire nw02405;
  wire nw02406;
  wire nw02407;
  wire nw02408;
  wire nw02409;
  wire nw02410;
  wire nw02411;
  wire nw02412;
  wire nw02413;
  wire nw02414;
  wire nw02415;
  wire nw02416;
  wire nw02417;
  wire nw02418;
  wire nw02419;
  wire nw02420;
  wire nw02421;
  wire nw02422;
  wire nw02423;
  wire nw02424;
  wire nw02425;
  wire nw02426;
  wire nw02427;
  wire nw02428;
  wire nw02429;
  wire nw02430;
  wire nw02431;
  wire nw02432;
  wire nw02433;
  wire nw02434;
  wire nw02435;
  wire nw02436;
  wire nw02437;
  wire nw02438;
  wire nw02439;
  wire nw02440;
  wire nw02441;
  wire nw02442;
  wire nw02443;
  wire nw02444;
  wire nw02445;
  wire nw02446;
  wire nw02447;
  wire nw02448;
  wire nw02449;
  wire nw02450;
  wire nw02451;
  wire nw02452;
  wire nw02453;
  wire nw02454;
  wire nw02455;
  wire nw02456;
  wire nw02457;
  wire nw02458;
  wire nw02459;
  wire nw02460;
  wire nw02461;
  wire nw02462;
  wire nw02463;
  wire nw02464;
  wire nw02465;
  wire nw02466;
  wire nw02467;
  wire nw02468;
  wire nw02469;
  wire nw02470;
  wire nw02471;
  wire nw02472;
  wire nw02473;
  wire nw02474;
  wire nw02475;
  wire nw02476;
  wire nw02477;
  wire nw02478;
  wire nw02479;
  wire nw02480;
  wire nw02481;
  wire nw02482;
  wire nw02483;
  wire nw02484;
  wire nw02485;
  wire nw02486;
  wire nw02487;
  wire nw02488;
  wire nw02489;
  wire nw02490;
  wire nw02491;
  wire nw02492;
  wire nw02493;
  wire nw02494;
  wire nw02495;
  wire nw02496;
  wire nw02497;
  wire nw02498;
  wire nw02499;
  wire nw02500;
  wire nw02501;
  wire nw02502;
  wire nw02503;
  wire nw02504;
  wire nw02505;
  wire nw02506;
  wire nw02507;
  wire nw02508;
  wire nw02509;
  wire nw02510;
  wire nw02511;
  wire nw02512;
  wire nw02513;
  wire nw02514;
  wire nw02515;
  wire nw02516;
  wire nw02517;
  wire nw02518;
  wire nw02519;
  wire nw02520;
  wire nw02521;
  wire nw02522;
  wire nw02523;
  wire nw02524;
  wire nw02525;
  wire nw02526;
  wire nw02527;
  wire nw02528;
  wire nw02529;
  wire nw02530;
  wire nw02531;
  wire nw02532;
  wire nw02533;
  wire nw02534;
  wire nw02535;
  wire nw02536;
  wire nw02537;
  wire nw02538;
  wire nw02539;
  wire nw02540;
  wire nw02541;
  wire nw02542;
  wire nw02543;
  wire nw02544;
  wire nw02545;
  wire nw02546;
  wire nw02547;
  wire nw02548;
  wire nw02549;
  wire nw02550;
  wire nw02551;
  wire nw02552;
  wire nw02553;
  wire nw02554;
  wire nw02555;
  wire nw02556;
  wire nw02557;
  wire nw02558;
  wire nw02559;
  wire nw02560;
  wire nw02561;
  wire nw02562;
  wire nw02563;
  wire nw02564;
  wire nw02565;
  wire nw02566;
  wire nw02567;
  wire nw02568;
  wire nw02569;
  wire nw02570;
  wire nw02571;
  wire nw02572;
  wire nw02573;
  wire nw02574;
  wire nw02575;
  wire nw02576;
  wire nw02577;
  wire nw02578;
  wire nw02579;
  wire nw02580;
  wire nw02581;
  wire nw02582;
  wire nw02583;
  wire nw02584;
  wire nw02585;
  wire nw02586;
  wire nw02587;
  wire nw02588;
  wire nw02589;
  wire nw02590;
  wire nw02591;
  wire nw02592;
  wire nw02593;
  wire nw02594;
  wire nw02595;
  wire nw02596;
  wire nw02597;
  wire nw02598;
  wire nw02599;
  wire nw02600;
  wire nw02601;
  wire nw02602;
  wire nw02603;
  wire nw02604;
  wire nw02605;
  wire nw02606;
  wire nw02607;
  wire nw02608;
  wire nw02609;
  wire nw02610;
  wire nw02611;
  wire nw02612;
  wire nw02613;
  wire nw02614;
  wire nw02615;
  wire nw02616;
  wire nw02617;
  wire nw02618;
  wire nw02619;
  wire nw02620;
  wire nw02621;
  wire nw02622;
  wire nw02623;
  wire nw02624;
  wire nw02625;
  wire nw02626;
  wire nw02627;
  wire nw02628;
  wire nw02629;
  wire nw02630;
  wire nw02631;
  wire nw02632;
  wire nw02633;
  wire nw02634;
  wire nw02635;
  wire nw02636;
  wire nw02637;
  wire nw02638;
  wire nw02639;
  wire nw02640;
  wire nw02641;
  wire nw02642;
  wire nw02643;
  wire nw02644;
  wire nw02645;
  wire nw02646;
  wire nw02647;
  wire nw02648;
  wire nw02649;
  wire nw02650;
  wire nw02651;
  wire nw02652;
  wire nw02653;
  wire nw02654;
  wire nw02655;
  wire nw02656;
  wire nw02657;
  wire nw02658;
  wire nw02659;
  wire nw02660;
  wire nw02661;
  wire nw02662;
  wire nw02663;
  wire nw02664;
  wire nw02665;
  wire nw02666;
  wire nw02667;
  wire nw02668;
  wire nw02669;
  wire nw02670;
  wire nw02671;
  wire nw02672;
  wire nw02673;
  wire nw02674;
  wire nw02675;
  wire nw02676;
  wire nw02677;
  wire nw02678;
  wire nw02679;
  wire nw02680;
  wire nw02681;
  wire nw02682;
  wire nw02683;
  wire nw02684;
  wire nw02685;
  wire nw02686;
  wire nw02687;
  wire nw02688;
  wire nw02689;
  wire nw02690;
  wire nw02691;
  wire nw02692;
  wire nw02693;
  wire nw02694;
  wire nw02695;
  wire nw02696;
  wire nw02697;
  wire nw02698;
  wire nw02699;
  wire nw02700;
  wire nw02701;
  wire nw02702;
  wire nw02703;
  wire nw02704;
  wire nw02705;
  wire nw02706;
  wire nw02707;
  wire nw02708;
  wire nw02709;
  wire nw02710;
  wire nw02711;
  wire nw02712;
  wire nw02713;
  wire nw02714;
  wire nw02715;
  wire nw02716;
  wire nw02717;
  wire nw02718;
  wire nw02719;
  wire nw02720;
  wire nw02721;
  wire nw02722;
  wire nw02723;
  wire nw02724;
  wire nw02725;
  wire nw02726;
  wire nw02727;
  wire nw02728;
  wire nw02729;
  wire nw02730;
  wire nw02731;
  wire nw02732;
  wire nw02733;
  wire nw02734;
  wire nw02735;
  wire nw02736;
  wire nw02737;
  wire nw02738;
  wire nw02739;
  wire nw02740;
  wire nw02741;
  wire nw02742;
  wire nw02743;
  wire nw02744;
  wire nw02745;
  wire nw02746;
  wire nw02747;
  wire nw02748;
  wire nw02749;
  wire nw02750;
  wire nw02751;
  wire nw02752;
  wire nw02753;
  wire nw02754;
  wire nw02755;
  wire nw02756;
  wire nw02757;
  wire nw02758;
  wire nw02759;
  wire nw02760;
  wire nw02761;
  wire nw02762;
  wire nw02763;
  wire nw02764;
  wire nw02765;
  wire nw02766;
  wire nw02767;
  wire nw02768;
  wire nw02769;
  wire nw02770;
  wire nw02771;
  wire nw02772;
  wire nw02773;
  wire nw02774;
  wire nw02775;
  wire nw02776;
  wire nw02777;
  wire nw02778;
  wire nw02779;
  wire nw02780;
  wire nw02781;
  wire nw02782;
  wire nw02783;
  wire nw02784;
  wire nw02785;
  wire nw02786;
  wire nw02787;
  wire nw02788;
  wire nw02789;
  wire nw02790;
  wire nw02791;
  wire nw02792;
  wire nw02793;
  wire nw02794;
  wire nw02795;
  wire nw02796;
  wire nw02797;
  wire nw02798;
  wire nw02799;
  wire nw02800;
  wire nw02801;
  wire nw02802;
  wire nw02803;
  wire nw02804;
  wire nw02805;
  wire nw02806;
  wire nw02807;
  wire nw02808;
  wire nw02809;
  wire nw02810;
  wire nw02811;
  wire nw02812;
  wire nw02813;
  wire nw02814;
  wire nw02815;
  wire nw02816;
  wire nw02817;
  wire nw02818;
  wire nw02819;
  wire nw02820;
  wire nw02821;
  wire nw02822;
  wire nw02823;
  wire nw02824;
  wire nw02825;
  wire nw02826;
  wire nw02827;
  wire nw02828;
  wire nw02829;
  wire nw02830;
  wire nw02831;
  wire nw02832;
  wire nw02833;
  wire nw02834;
  wire nw02835;
  wire nw02836;
  wire nw02837;
  wire nw02838;
  wire nw02839;
  wire nw02840;
  wire nw02841;
  wire nw02842;
  wire nw02843;
  wire nw02844;
  wire nw02845;
  wire nw02846;
  wire nw02847;
  wire nw02848;
  wire nw02849;
  wire nw02850;
  wire nw02851;
  wire nw02852;
  wire nw02853;
  wire nw02854;
  wire nw02855;
  wire nw02856;
  wire nw02857;
  wire nw02858;
  wire nw02859;
  wire nw02860;
  wire nw02861;
  wire nw02862;
  wire nw02863;
  wire nw02864;
  wire nw02865;
  wire nw02866;
  wire nw02867;
  wire nw02868;
  wire nw02869;
  wire nw02870;
  wire nw02871;
  wire nw02872;
  wire nw02873;
  wire nw02874;
  wire nw02875;
  wire nw02876;
  wire nw02877;
  wire nw02878;
  wire nw02879;
  wire nw02880;
  wire nw02881;
  wire nw02882;
  wire nw02883;
  wire nw02884;
  wire nw02885;
  wire nw02886;
  wire nw02887;
  wire nw02888;
  wire nw02889;
  wire nw02890;
  wire nw02891;
  wire nw02892;
  wire nw02893;
  wire nw02894;
  wire nw02895;
  wire nw02896;
  wire nw02897;
  wire nw02898;
  wire nw02899;
  wire nw02900;
  wire nw02901;
  wire nw02902;
  wire nw02903;
  wire nw02904;
  wire nw02905;
  wire nw02906;
  wire nw02907;
  wire nw02908;
  wire nw02909;
  wire nw02910;
  wire nw02911;
  wire nw02912;
  wire nw02913;
  wire nw02914;
  wire nw02915;
  wire nw02916;
  wire nw02917;
  wire nw02918;
  wire nw02919;
  wire nw02920;
  wire nw02921;
  wire nw02922;
  wire nw02923;
  wire nw02924;
  wire nw02925;
  wire nw02926;
  wire nw02927;
  wire nw02928;
  wire nw02929;
  wire nw02930;
  wire nw02931;
  wire nw02932;
  wire nw02933;
  wire nw02934;
  wire nw02935;
  wire nw02936;
  wire nw02937;
  wire nw02938;
  wire nw02939;
  wire nw02940;
  wire nw02941;
  wire nw02942;
  wire nw02943;
  wire nw02944;
  wire nw02945;
  wire nw02946;
  wire nw02947;
  wire nw02948;
  wire nw02949;
  wire nw02950;
  wire nw02951;
  wire nw02952;
  wire nw02953;
  wire nw02954;
  wire nw02955;
  wire nw02956;
  wire nw02957;
  wire nw02958;
  wire nw02959;
  wire nw02960;
  wire nw02961;
  wire nw02962;
  wire nw02963;
  wire nw02964;
  wire nw02965;
  wire nw02966;
  wire nw02967;
  wire nw02968;
  wire nw02969;
  wire nw02970;
  wire nw02971;
  wire nw02972;
  wire nw02973;
  wire nw02974;
  wire nw02975;
  wire nw02976;
  wire nw02977;
  wire nw02978;
  wire nw02979;
  wire nw02980;
  wire nw02981;
  wire nw02982;
  wire nw02983;
  wire nw02984;
  wire nw02985;
  wire nw02986;
  wire nw02987;
  wire nw02988;
  wire nw02989;
  wire nw02990;
  wire nw02991;
  wire nw02992;
  wire nw02993;
  wire nw02994;
  wire nw02995;
  wire nw02996;
  wire nw02997;
  wire nw02998;
  wire nw02999;
  wire nw03000;
  wire nw03001;
  wire nw03002;
  wire nw03003;
  wire nw03004;
  wire nw03005;
  wire nw03006;
  wire nw03007;
  wire nw03008;
  wire nw03009;
  wire nw03010;
  wire nw03011;
  wire nw03012;
  wire nw03013;
  wire nw03014;
  wire nw03015;
  wire nw03016;
  wire nw03017;
  wire nw03018;
  wire nw03019;
  wire nw03020;
  wire nw03021;
  wire nw03022;
  wire nw03023;
  wire nw03024;
  wire nw03025;
  wire nw03026;
  wire nw03027;
  wire nw03028;
  wire nw03029;
  wire nw03030;
  wire nw03031;
  wire nw03032;
  wire nw03033;
  wire nw03034;
  wire nw03035;
  wire nw03036;
  wire nw03037;
  wire nw03038;
  wire nw03039;
  wire nw03040;
  wire nw03041;
  wire nw03042;
  wire nw03043;
  wire nw03044;
  wire nw03045;
  wire nw03046;
  wire nw03047;
  wire nw03048;
  wire nw03049;
  wire nw03050;
  wire nw03051;
  wire nw03052;
  wire nw03053;
  wire nw03054;
  wire nw03055;
  wire nw03056;
  wire nw03057;
  wire nw03058;
  wire nw03059;
  wire nw03060;
  wire nw03061;
  wire nw03062;
  wire nw03063;
  wire nw03064;
  wire nw03065;
  wire nw03066;
  wire nw03067;
  wire nw03068;
  wire nw03069;
  wire nw03070;
  wire nw03071;
  wire nw03072;
  wire nw03073;
  wire nw03074;
  wire nw03075;
  wire nw03076;
  wire nw03077;
  wire nw03078;
  wire nw03079;
  wire nw03080;
  wire nw03081;
  wire nw03082;
  wire nw03083;
  wire nw03084;
  wire nw03085;
  wire nw03086;
  wire nw03087;
  wire nw03088;
  wire nw03089;
  wire nw03090;
  wire nw03091;
  wire nw03092;
  wire nw03093;
  wire nw03094;
  wire nw03095;
  wire nw03096;
  wire nw03097;
  wire nw03098;
  wire nw03099;
  wire nw03100;
  wire nw03101;
  wire nw03102;
  wire nw03103;
  wire nw03104;
  wire nw03105;
  wire nw03106;
  wire nw03107;
  wire nw03108;
  wire nw03109;
  wire nw03110;
  wire nw03111;
  wire nw03112;
  wire nw03113;
  wire nw03114;
  wire nw03115;
  wire nw03116;
  wire nw03117;
  wire nw03118;
  wire nw03119;
  wire nw03120;
  wire nw03121;
  wire nw03122;
  wire nw03123;
  wire nw03124;
  wire nw03125;
  wire nw03126;
  wire nw03127;
  wire nw03128;
  wire nw03129;
  wire nw03130;
  wire nw03131;
  wire nw03132;
  wire nw03133;
  wire nw03134;
  wire nw03135;
  wire nw03136;
  wire nw03137;
  wire nw03138;
  wire nw03139;
  wire nw03140;
  wire nw03141;
  wire nw03142;
  wire nw03143;
  wire nw03144;
  wire nw03145;
  wire nw03146;
  wire nw03147;
  wire nw03148;
  wire nw03149;
  wire nw03150;
  wire nw03151;
  wire nw03152;
  wire nw03153;
  wire nw03154;
  wire nw03155;
  wire nw03156;
  wire nw03157;
  wire nw03158;
  wire nw03159;
  wire nw03160;
  wire nw03161;
  wire nw03162;
  wire nw03163;
  wire nw03164;
  wire nw03165;
  wire nw03166;
  wire nw03167;
  wire nw03168;
  wire nw03169;
  wire nw03170;
  wire nw03171;
  wire nw03172;
  wire nw03173;
  wire nw03174;
  wire nw03175;
  wire nw03176;
  wire nw03177;
  wire nw03178;
  wire nw03179;
  wire nw03180;
  wire nw03181;
  wire nw03182;
  wire nw03183;
  wire nw03184;
  wire nw03185;
  wire nw03186;
  wire nw03187;
  wire nw03188;
  wire nw03189;
  wire nw03190;
  wire nw03191;
  wire nw03192;
  wire nw03193;
  wire nw03194;
  wire nw03195;
  wire nw03196;
  wire nw03197;
  wire nw03198;
  wire nw03199;
  wire nw03200;
  wire nw03201;
  wire nw03202;
  wire nw03203;
  wire nw03204;
  wire nw03205;
  wire nw03206;
  wire nw03207;
  wire nw03208;
  wire nw03209;
  wire nw03210;
  wire nw03211;
  wire nw03212;
  wire nw03213;
  wire nw03214;
  wire nw03215;
  wire nw03216;
  wire nw03217;
  wire nw03218;
  wire nw03219;
  wire nw03220;
  wire nw03221;
  wire nw03222;
  wire nw03223;
  wire nw03224;
  wire nw03225;
  wire nw03226;
  wire nw03227;
  wire nw03228;
  wire nw03229;
  wire nw03230;
  wire nw03231;
  wire nw03232;
  wire nw03233;
  wire nw03234;
  wire nw03235;
  wire nw03236;
  wire nw03237;
  wire nw03238;
  wire nw03239;
  wire nw03240;
  wire nw03241;
  wire nw03242;
  wire nw03243;
  wire nw03244;
  wire nw03245;
  wire nw03246;
  wire nw03247;
  wire nw03248;
  wire nw03249;
  wire nw03250;
  wire nw03251;
  wire nw03252;
  wire nw03253;
  wire nw03254;
  wire nw03255;
  wire nw03256;
  wire nw03257;
  wire nw03258;
  wire nw03259;
  wire nw03260;
  wire nw03261;
  wire nw03262;
  wire nw03263;
  wire nw03264;
  wire nw03265;
  wire nw03266;
  wire nw03267;
  wire nw03268;
  wire nw03269;
  wire nw03270;
  wire nw03271;
  wire nw03272;
  wire nw03273;
  wire nw03274;
  wire nw03275;
  wire nw03276;
  wire nw03277;
  wire nw03278;
  wire nw03279;
  wire nw03280;
  wire nw03281;
  wire nw03282;
  wire nw03283;
  wire nw03284;
  wire nw03285;
  wire nw03286;
  wire nw03287;
  wire nw03288;
  wire nw03289;
  wire nw03290;
  wire nw03291;
  wire nw03292;
  wire nw03293;
  wire nw03294;
  wire nw03295;
  wire nw03296;
  wire nw03297;
  wire nw03298;
  wire nw03299;
  wire nw03300;
  wire nw03301;
  wire nw03302;
  wire nw03303;
  wire nw03304;
  wire nw03305;
  wire nw03306;
  wire nw03307;
  wire nw03308;
  wire nw03309;
  wire nw03310;
  wire nw03311;
  wire nw03312;
  wire nw03313;
  wire nw03314;
  wire nw03315;
  wire nw03316;
  wire nw03317;
  wire nw03318;
  wire nw03319;
  wire nw03320;
  wire nw03321;
  wire nw03322;
  wire nw03323;
  wire nw03324;
  wire nw03325;
  wire nw03326;
  wire nw03327;
  wire nw03328;
  wire nw03329;
  wire nw03330;
  wire nw03331;
  wire nw03332;
  wire nw03333;
  wire nw03334;
  wire nw03335;
  wire nw03336;
  wire nw03337;
  wire nw03338;
  wire nw03339;
  wire nw03340;
  wire nw03341;
  wire nw03342;
  wire nw03343;
  wire nw03344;
  wire nw03345;
  wire nw03346;
  wire nw03347;
  wire nw03348;
  wire nw03349;
  wire nw03350;
  wire nw03351;
  wire nw03352;
  wire nw03353;
  wire nw03354;
  wire nw03355;
  wire nw03356;
  wire nw03357;
  wire nw03358;
  wire nw03359;
  wire nw03360;
  wire nw03361;
  wire nw03362;
  wire nw03363;
  wire nw03364;
  wire nw03365;
  wire nw03366;
  wire nw03367;
  wire nw03368;
  wire nw03369;
  wire nw03370;
  wire nw03371;
  wire nw03372;
  wire nw03373;
  wire nw03374;
  wire nw03375;
  wire nw03376;
  wire nw03377;
  wire nw03378;
  wire nw03379;
  wire nw03380;
  wire nw03381;
  wire nw03382;
  wire nw03383;
  wire nw03384;
  wire nw03385;
  wire nw03386;
  wire nw03387;
  wire nw03388;
  wire nw03389;
  wire nw03390;
  wire nw03391;
  wire nw03392;
  wire nw03393;
  wire nw03394;
  wire nw03395;
  wire nw03396;
  wire nw03397;
  wire nw03398;
  wire nw03399;
  wire nw03400;
  wire nw03401;
  wire nw03402;
  wire nw03403;
  wire nw03404;
  wire nw03405;
  wire nw03406;
  wire nw03407;
  wire nw03408;
  wire nw03409;
  wire nw03410;
  wire nw03411;
  wire nw03412;
  wire nw03413;
  wire nw03414;
  wire nw03415;
  wire nw03416;
  wire nw03417;
  wire nw03418;
  wire nw03419;
  wire nw03420;
  wire nw03421;
  wire nw03422;
  wire nw03423;
  wire nw03424;
  wire nw03425;
  wire nw03426;
  wire nw03427;
  wire nw03428;
  wire nw03429;
  wire nw03430;
  wire nw03431;
  wire nw03432;
  wire nw03433;
  wire nw03434;
  wire nw03435;
  wire nw03436;
  wire nw03437;
  wire nw03438;
  wire nw03439;
  wire nw03440;
  wire nw03441;
  wire nw03442;
  wire nw03443;
  wire nw03444;
  wire nw03445;
  wire nw03446;
  wire nw03447;
  wire nw03448;
  wire nw03449;
  wire nw03450;
  wire nw03451;
  wire nw03452;
  wire nw03453;
  wire nw03454;
  wire nw03455;
  wire nw03456;
  wire nw03457;
  wire nw03458;
  wire nw03459;
  wire nw03460;
  wire nw03461;
  wire nw03462;
  wire nw03463;
  wire nw03464;
  wire nw03465;
  wire nw03466;
  wire nw03467;
  wire nw03468;
  wire nw03469;
  wire nw03470;
  wire nw03471;
  wire nw03472;
  wire nw03473;
  wire nw03474;
  wire nw03475;
  wire nw03476;
  wire nw03477;
  wire nw03478;
  wire nw03479;
  wire nw03480;
  wire nw03481;
  wire nw03482;
  wire nw03483;
  wire nw03484;
  wire nw03485;
  wire nw03486;
  wire nw03487;
  wire nw03488;
  wire nw03489;
  wire nw03490;
  wire nw03491;
  wire nw03492;
  wire nw03493;
  wire nw03494;
  wire nw03495;
  wire nw03496;
  wire nw03497;
  wire nw03498;
  wire nw03499;
  wire nw03500;
  wire nw03501;
  wire nw03502;
  wire nw03503;
  wire nw03504;
  wire nw03505;
  wire nw03506;
  wire nw03507;
  wire nw03508;
  wire nw03509;
  wire nw03510;
  wire nw03511;
  wire nw03512;
  wire nw03513;
  wire nw03514;
  wire nw03515;
  wire nw03516;
  wire nw03517;
  wire nw03518;
  wire nw03519;
  wire nw03520;
  wire nw03521;
  wire nw03522;
  wire nw03523;
  wire nw03524;
  wire nw03525;
  wire nw03526;
  wire nw03527;
  wire nw03528;
  wire nw03529;
  wire nw03530;
  wire nw03531;
  wire nw03532;
  wire nw03533;
  wire nw03534;
  wire nw03535;
  wire nw03536;
  wire nw03537;
  wire nw03538;
  wire nw03539;
  wire nw03540;
  wire nw03541;
  wire nw03542;
  wire nw03543;
  wire nw03544;
  wire nw03545;
  wire nw03546;
  wire nw03547;
  wire nw03548;
  wire nw03549;
  wire nw03550;
  wire nw03551;
  wire nw03552;
  wire nw03553;
  wire nw03554;
  wire nw03555;
  wire nw03556;
  wire nw03557;
  wire nw03558;
  wire nw03559;
  wire nw03560;
  wire nw03561;
  wire nw03562;
  wire nw03563;
  wire nw03564;
  wire nw03565;
  wire nw03566;
  wire nw03567;
  wire nw03568;
  wire nw03569;
  wire nw03570;
  wire nw03571;
  wire nw03572;
  wire nw03573;
  wire nw03574;
  wire nw03575;
  wire nw03576;
  wire nw03577;
  wire nw03578;
  wire nw03579;
  wire nw03580;
  wire nw03581;
  wire nw03582;
  wire nw03583;
  wire nw03584;
  wire nw03585;
  wire nw03586;
  wire nw03587;
  wire nw03588;
  wire nw03589;
  wire nw03590;
  wire nw03591;
  wire nw03592;
  wire nw03593;
  wire nw03594;
  wire nw03595;
  wire nw03596;
  wire nw03597;
  wire nw03598;
  wire nw03599;
  wire nw03600;
  wire nw03601;
  wire nw03602;
  wire nw03603;
  wire nw03604;
  wire nw03605;
  wire nw03606;
  wire nw03607;
  wire nw03608;
  wire nw03609;
  wire nw03610;
  wire nw03611;
  wire nw03612;
  wire nw03613;
  wire nw03614;
  wire nw03615;
  wire nw03616;
  wire nw03617;
  wire nw03618;
  wire nw03619;
  wire nw03620;
  wire nw03621;
  wire nw03622;
  wire nw03623;
  wire nw03624;
  wire nw03625;
  wire nw03626;
  wire nw03627;
  wire nw03628;
  wire nw03629;
  wire nw03630;
  wire nw03631;
  wire nw03632;
  wire nw03633;
  wire nw03634;
  wire nw03635;
  wire nw03636;
  wire nw03637;
  wire nw03638;
  wire nw03639;
  wire nw03640;
  wire nw03641;
  wire nw03642;
  wire nw03643;
  wire nw03644;
  wire nw03645;
  wire nw03646;
  wire nw03647;
  wire nw03648;
  wire nw03649;
  wire nw03650;
  wire nw03651;
  wire nw03652;
  wire nw03653;
  wire nw03654;
  wire nw03655;
  wire nw03656;
  wire nw03657;
  wire nw03658;
  wire nw03659;
  wire nw03660;
  wire nw03661;
  wire nw03662;
  wire nw03663;
  wire nw03664;
  wire nw03665;
  wire nw03666;
  wire nw03667;
  wire nw03668;
  wire nw03669;
  wire nw03670;
  wire nw03671;
  wire nw03672;
  wire nw03673;
  wire nw03674;
  wire nw03675;
  wire nw03676;
  wire nw03677;
  wire nw03678;
  wire nw03679;
  wire nw03680;
  wire nw03681;
  wire nw03682;
  wire nw03683;
  wire nw03684;
  wire nw03685;
  wire nw03686;
  wire nw03687;
  wire nw03688;
  wire nw03689;
  wire nw03690;
  wire nw03691;
  wire nw03692;
  wire nw03693;
  wire nw03694;
  wire nw03695;
  wire nw03696;
  wire nw03697;
  wire nw03698;
  wire nw03699;
  wire nw03700;
  wire nw03701;
  wire nw03702;
  wire nw03703;
  wire nw03704;
  wire nw03705;
  wire nw03706;
  wire nw03707;
  wire nw03708;
  wire nw03709;
  wire nw03710;
  wire nw03711;
  wire nw03712;
  wire nw03713;
  wire nw03714;
  wire nw03715;
  wire nw03716;
  wire nw03717;
  wire nw03718;
  wire nw03719;
  wire nw03720;
  wire nw03721;
  wire nw03722;
  wire nw03723;
  wire nw03724;
  wire nw03725;
  wire nw03726;
  wire nw03727;
  wire nw03728;
  wire nw03729;
  wire nw03730;
  wire nw03731;
  wire nw03732;
  wire nw03733;
  wire nw03734;
  wire nw03735;
  wire nw03736;
  wire nw03737;
  wire nw03738;
  wire nw03739;
  wire nw03740;
  wire nw03741;
  wire nw03742;
  wire nw03743;
  wire nw03744;
  wire nw03745;
  wire nw03746;
  wire nw03747;
  wire nw03748;
  wire nw03749;
  wire nw03750;
  wire nw03751;
  wire nw03752;
  wire nw03753;
  wire nw03754;
  wire nw03755;
  wire nw03756;
  wire nw03757;
  wire nw03758;
  wire nw03759;
  wire nw03760;
  wire nw03761;
  wire nw03762;
  wire nw03763;
  wire nw03764;
  wire nw03765;
  wire nw03766;
  wire nw03767;
  wire nw03768;
  wire nw03769;
  wire nw03770;
  wire nw03771;
  wire nw03772;
  wire nw03773;
  wire nw03774;
  wire nw03775;
  wire nw03776;
  wire nw03777;
  wire nw03778;
  wire nw03779;
  wire nw03780;
  wire nw03781;
  wire nw03782;
  wire nw03783;
  wire nw03784;
  wire nw03785;
  wire nw03786;
  wire nw03787;
  wire nw03788;
  wire nw03789;
  wire nw03790;
  wire nw03791;
  wire nw03792;
  wire nw03793;
  wire nw03794;
  wire nw03795;
  wire nw03796;
  wire nw03797;
  wire nw03798;
  wire nw03799;
  wire nw03800;
  wire nw03801;
  wire nw03802;
  wire nw03803;
  wire nw03804;
  wire nw03805;
  wire nw03806;
  wire nw03807;
  wire nw03808;
  wire nw03809;
  wire nw03810;
  wire nw03811;
  wire nw03812;
  wire nw03813;
  wire nw03814;
  wire nw03815;
  wire nw03816;
  wire nw03817;
  wire nw03818;
  wire nw03819;
  wire nw03820;
  wire nw03821;
  wire nw03822;
  wire nw03823;
  wire nw03824;
  wire nw03825;
  wire nw03826;
  wire nw03827;
  wire nw03828;
  wire nw03829;
  wire nw03830;
  wire nw03831;
  wire nw03832;
  wire nw03833;
  wire nw03834;
  wire nw03835;
  wire nw03836;
  wire nw03837;
  wire nw03838;
  wire nw03839;
  wire nw03840;
  wire nw03841;
  wire nw03842;
  wire nw03843;
  wire nw03844;
  wire nw03845;
  wire nw03846;
  wire nw03847;
  wire nw03848;
  wire nw03849;
  wire nw03850;
  wire nw03851;
  wire nw03852;
  wire nw03853;
  wire nw03854;
  wire nw03855;
  wire nw03856;
  wire nw03857;
  wire nw03858;
  wire nw03859;
  wire nw03860;
  wire nw03861;
  wire nw03862;
  wire nw03863;
  wire nw03864;
  wire nw03865;
  wire nw03866;
  wire nw03867;
  wire nw03868;
  wire nw03869;
  wire nw03870;
  wire nw03871;
  wire nw03872;
  wire nw03873;
  wire nw03874;
  wire nw03875;
  wire nw03876;
  wire nw03877;
  wire nw03878;
  wire nw03879;
  wire nw03880;
  wire nw03881;
  wire nw03882;
  wire nw03883;
  wire nw03884;
  wire nw03885;
  wire nw03886;
  wire nw03887;
  wire nw03888;
  wire nw03889;
  wire nw03890;
  wire nw03891;
  wire nw03892;
  wire nw03893;
  wire nw03894;
  wire nw03895;
  wire nw03896;
  wire nw03897;
  wire nw03898;
  wire nw03899;
  wire nw03900;
  wire nw03901;
  wire nw03902;
  wire nw03903;
  wire nw03904;
  wire nw03905;
  wire nw03906;
  wire nw03907;
  wire nw03908;
  wire nw03909;
  wire nw03910;
  wire nw03911;
  wire nw03912;
  wire nw03913;
  wire nw03914;
  wire nw03915;
  wire nw03916;
  wire nw03917;
  wire nw03918;
  wire nw03919;
  wire nw03920;
  wire nw03921;
  wire nw03922;
  wire nw03923;
  wire nw03924;
  wire nw03925;
  wire nw03926;
  wire nw03927;
  wire nw03928;
  wire nw03929;
  wire nw03930;
  wire nw03931;
  wire nw03932;
  wire nw03933;
  wire nw03934;
  wire nw03935;
  wire nw03936;
  wire nw03937;
  wire nw03938;
  wire nw03939;
  wire nw03940;
  wire nw03941;
  wire nw03942;
  wire nw03943;
  wire nw03944;
  wire nw03945;
  wire nw03946;
  wire nw03947;
  wire nw03948;
  wire nw03949;
  wire nw03950;
  wire nw03951;
  wire nw03952;
  wire nw03953;
  wire nw03954;
  wire nw03955;
  wire nw03956;
  wire nw03957;
  wire nw03958;
  wire nw03959;
  wire nw03960;
  wire nw03961;
  wire nw03962;
  wire nw03963;
  wire nw03964;
  wire nw03965;
  wire nw03966;
  wire nw03967;
  wire nw03968;
  wire nw03969;
  wire nw03970;
  wire nw03971;
  wire nw03972;
  wire nw03973;
  wire nw03974;
  wire nw03975;
  wire nw03976;
  wire nw03977;
  wire nw03978;
  wire nw03979;
  wire nw03980;
  wire nw03981;
  wire nw03982;
  wire nw03983;
  wire nw03984;
  wire nw03985;
  wire nw03986;
  wire nw03987;
  wire nw03988;
  wire nw03989;
  wire nw03990;
  wire nw03991;
  wire nw03992;
  wire nw03993;
  wire nw03994;
  wire nw03995;
  wire nw03996;
  wire nw03997;
  wire nw03998;
  wire nw03999;
  wire nw04000;
  wire nw04001;
  wire nw04002;
  wire nw04003;
  wire nw04004;
  wire nw04005;
  wire nw04006;
  wire nw04007;
  wire nw04008;
  wire nw04009;
  wire nw04010;
  wire nw04011;
  wire nw04012;
  wire nw04013;
  wire nw04014;
  wire nw04015;
  wire nw04016;
  wire nw04017;
  wire nw04018;
  wire nw04019;
  wire nw04020;
  wire nw04021;
  wire nw04022;
  wire nw04023;
  wire nw04024;
  wire nw04025;
  wire nw04026;
  wire nw04027;
  wire nw04028;
  wire nw04029;
  wire nw04030;
  wire nw04031;
  wire nw04032;
  wire nw04033;
  wire nw04034;
  wire nw04035;
  wire nw04036;
  wire nw04037;
  wire nw04038;
  wire nw04039;
  wire nw04040;
  wire nw04041;
  wire nw04042;
  wire nw04043;
  wire nw04044;
  wire nw04045;
  wire nw04046;
  wire nw04047;
  wire nw04048;
  wire nw04049;
  wire nw04050;
  wire nw04051;
  wire nw04052;
  wire nw04053;
  wire nw04054;
  wire nw04055;
  wire nw04056;
  wire nw04057;
  wire nw04058;
  wire nw04059;
  wire nw04060;
  wire nw04061;
  wire nw04062;
  wire nw04063;
  wire nw04064;
  wire nw04065;
  wire nw04066;
  wire nw04067;
  wire nw04068;
  wire nw04069;
  wire nw04070;
  wire nw04071;
  wire nw04072;
  wire nw04073;
  wire nw04074;
  wire nw04075;
  wire nw04076;
  wire nw04077;
  wire nw04078;
  wire nw04079;
  wire nw04080;
  wire nw04081;
  wire nw04082;
  wire nw04083;
  wire nw04084;
  wire nw04085;
  wire nw04086;
  wire nw04087;
  wire nw04088;
  wire nw04089;
  wire nw04090;
  wire nw04091;
  wire nw04092;
  wire nw04093;
  wire nw04094;
  wire nw04095;
  wire nw04096;
  wire nw04097;
  wire nw04098;
  wire nw04099;
  wire nw04100;
  wire nw04101;
  wire nw04102;
  wire nw04103;
  wire nw04104;
  wire nw04105;
  wire nw04106;
  wire nw04107;
  wire nw04108;
  wire nw04109;
  wire nw04110;
  wire nw04111;
  wire nw04112;
  wire nw04113;
  wire nw04114;
  wire nw04115;
  wire nw04116;
  wire nw04117;
  wire nw04118;
  wire nw04119;
  wire nw04120;
  wire nw04121;
  wire nw04122;
  wire nw04123;
  wire nw04124;
  wire nw04125;
  wire nw04126;
  wire nw04127;
  wire nw04128;
  wire nw04129;
  wire nw04130;
  wire nw04131;
  wire nw04132;
  wire nw04133;
  wire nw04134;
  wire nw04135;
  wire nw04136;
  wire nw04137;
  wire nw04138;
  wire nw04139;
  wire nw04140;
  wire nw04141;
  wire nw04142;
  wire nw04143;
  wire nw04144;
  wire nw04145;
  wire nw04146;
  wire nw04147;
  wire nw04148;
  wire nw04149;
  wire nw04150;
  wire nw04151;
  wire nw04152;
  wire nw04153;
  wire nw04154;
  wire nw04155;
  wire nw04156;
  wire nw04157;
  wire nw04158;
  wire nw04159;
  wire nw04160;
  wire nw04161;
  wire nw04162;
  wire nw04163;
  wire nw04164;
  wire nw04165;
  wire nw04166;
  wire nw04167;
  wire nw04168;
  wire nw04169;
  wire nw04170;
  wire nw04171;
  wire nw04172;
  wire nw04173;
  wire nw04174;
  wire nw04175;
  wire nw04176;
  wire nw04177;
  wire nw04178;
  wire nw04179;
  wire nw04180;
  wire nw04181;
  wire nw04182;
  wire nw04183;
  wire nw04184;
  wire nw04185;
  wire nw04186;
  wire nw04187;
  wire nw04188;
  wire nw04189;
  wire nw04190;
  wire nw04191;
  wire nw04192;
  wire nw04193;
  wire nw04194;
  wire nw04195;
  wire nw04196;
  wire nw04197;
  wire nw04198;
  wire nw04199;
  wire nw04200;
  wire nw04201;
  wire nw04202;
  wire nw04203;
  wire nw04204;
  wire nw04205;
  wire nw04206;
  wire nw04207;
  wire nw04208;
  wire nw04209;
  wire nw04210;
  wire nw04211;
  wire nw04212;
  wire nw04213;
  wire nw04214;
  wire nw04215;
  wire nw04216;
  wire nw04217;
  wire nw04218;
  wire nw04219;
  wire nw04220;
  wire nw04221;
  wire nw04222;
  wire nw04223;
  wire nw04224;
  wire nw04225;
  wire nw04226;
  wire nw04227;
  wire nw04228;
  wire nw04229;
  wire nw04230;
  wire nw04231;
  wire nw04232;
  wire nw04233;
  wire nw04234;
  wire nw04235;
  wire nw04236;
  wire nw04237;
  wire nw04238;
  wire nw04239;
  wire nw04240;
  wire nw04241;
  wire nw04242;
  wire nw04243;
  wire nw04244;
  wire nw04245;
  wire nw04246;
  wire nw04247;
  wire nw04248;
  wire nw04249;
  wire nw04250;
  wire nw04251;
  wire nw04252;
  wire nw04253;
  wire nw04254;
  wire nw04255;
  wire nw04256;
  wire nw04257;
  wire nw04258;
  wire nw04259;
  wire nw04260;
  wire nw04261;
  wire nw04262;
  wire nw04263;
  wire nw04264;
  wire nw04265;
  wire nw04266;
  wire nw04267;
  wire nw04268;
  wire nw04269;
  wire nw04270;
  wire nw04271;
  wire nw04272;
  wire nw04273;
  wire nw04274;
  wire nw04275;
  wire nw04276;
  wire nw04277;
  wire nw04278;
  wire nw04279;
  wire nw04280;
  wire nw04281;
  wire nw04282;
  wire nw04283;
  wire nw04284;
  wire nw04285;
  wire nw04286;
  wire nw04287;
  wire nw04288;
  wire nw04289;
  wire nw04290;
  wire nw04291;
  wire nw04292;
  wire nw04293;
  wire nw04294;
  wire nw04295;
  wire nw04296;
  wire nw04297;
  wire nw04298;
  wire nw04299;
  wire nw04300;
  wire nw04301;
  wire nw04302;
  wire nw04303;
  wire nw04304;
  wire nw04305;
  wire nw04306;
  wire nw04307;
  wire nw04308;
  wire nw04309;
  wire nw04310;
  wire nw04311;
  wire nw04312;
  wire nw04313;
  wire nw04314;
  wire nw04315;
  wire nw04316;
  wire nw04317;
  wire nw04318;
  wire nw04319;
  wire nw04320;
  wire nw04321;
  wire nw04322;
  wire nw04323;
  wire nw04324;
  wire nw04325;
  wire nw04326;
  wire nw04327;
  wire nw04328;
  wire nw04329;
  wire nw04330;
  wire nw04331;
  wire nw04332;
  wire nw04333;
  wire nw04334;
  wire nw04335;
  wire nw04336;
  wire nw04337;
  wire nw04338;
  wire nw04339;
  wire nw04340;
  wire nw04341;
  wire nw04342;
  wire nw04343;
  wire nw04344;
  wire nw04345;
  wire nw04346;
  wire nw04347;
  wire nw04348;
  wire nw04349;
  wire nw04350;
  wire nw04351;
  wire nw04352;
  wire nw04353;
  wire nw04354;
  wire nw04355;
  wire nw04356;
  wire nw04357;
  wire nw04358;
  wire nw04359;
  wire nw04360;
  wire nw04361;
  wire nw04362;
  wire nw04363;
  wire nw04364;
  wire nw04365;
  wire nw04366;
  wire nw04367;
  wire nw04368;
  wire nw04369;
  wire nw04370;
  wire nw04371;
  wire nw04372;
  wire nw04373;
  wire nw04374;
  wire nw04375;
  wire nw04376;
  wire nw04377;
  wire nw04378;
  wire nw04379;
  wire nw04380;
  wire nw04381;
  wire nw04382;
  wire nw04383;
  wire nw04384;
  wire nw04385;
  wire nw04386;
  wire nw04387;
  wire nw04388;
  wire nw04389;
  wire nw04390;
  wire nw04391;
  wire nw04392;
  wire nw04393;
  wire nw04394;
  wire nw04395;
  wire nw04396;
  wire nw04397;
  wire nw04398;
  wire nw04399;
  wire nw04400;
  wire nw04401;
  wire nw04402;
  wire nw04403;
  wire nw04404;
  wire nw04405;
  wire nw04406;
  wire nw04407;
  wire nw04408;
  wire nw04409;
  wire nw04410;
  wire nw04411;
  wire nw04412;
  wire nw04413;
  wire nw04414;
  wire nw04415;
  wire nw04416;
  wire nw04417;
  wire nw04418;
  wire nw04419;
  wire nw04420;
  wire nw04421;
  wire nw04422;
  wire nw04423;
  wire nw04424;
  wire nw04425;
  wire nw04426;
  wire nw04427;
  wire nw04428;
  wire nw04429;
  wire nw04430;
  wire nw04431;
  wire nw04432;
  wire nw04433;
  wire nw04434;
  wire nw04435;
  wire nw04436;
  wire nw04437;
  wire nw04438;
  wire nw04439;
  wire nw04440;
  wire nw04441;
  wire nw04442;
  wire nw04443;
  wire nw04444;
  wire nw04445;
  wire nw04446;
  wire nw04447;
  wire nw04448;
  wire nw04449;
  wire nw04450;
  wire nw04451;
  wire nw04452;
  wire nw04453;
  wire nw04454;
  wire nw04455;
  wire nw04456;
  wire nw04457;
  wire nw04458;
  wire nw04459;
  wire nw04460;
  wire nw04461;
  wire nw04462;
  wire nw04463;
  wire nw04464;
  wire nw04465;
  wire nw04466;
  wire nw04467;
  wire nw04468;
  wire nw04469;
  wire nw04470;
  wire nw04471;
  wire nw04472;
  wire nw04473;
  wire nw04474;
  wire nw04475;
  wire nw04476;
  wire nw04477;
  wire nw04478;
  wire nw04479;
  wire nw04480;
  wire nw04481;
  wire nw04482;
  wire nw04483;
  wire nw04484;
  wire nw04485;
  wire nw04486;
  wire nw04487;
  wire nw04488;
  wire nw04489;
  wire nw04490;
  wire nw04491;
  wire nw04492;
  wire nw04493;
  wire nw04494;
  wire nw04495;
  wire nw04496;
  wire nw04497;
  wire nw04498;
  wire nw04499;
  wire nw04500;
  wire nw04501;
  wire nw04502;
  wire nw04503;
  wire nw04504;
  wire nw04505;
  wire nw04506;
  wire nw04507;
  wire nw04508;
  wire nw04509;
  wire nw04510;
  wire nw04511;
  wire nw04512;
  wire nw04513;
  wire nw04514;
  wire nw04515;
  wire nw04516;
  wire nw04517;
  wire nw04518;
  wire nw04519;
  wire nw04520;
  wire nw04521;
  wire nw04522;
  wire nw04523;
  wire nw04524;
  wire nw04525;
  wire nw04526;
  wire nw04527;
  wire nw04528;
  wire nw04529;
  wire nw04530;
  wire nw04531;
  wire nw04532;
  wire nw04533;
  wire nw04534;
  wire nw04535;
  wire nw04536;
  wire nw04537;
  wire nw04538;
  wire nw04539;
  wire nw04540;
  wire nw04541;
  wire nw04542;
  wire nw04543;
  wire nw04544;
  wire nw04545;
  wire nw04546;
  wire nw04547;
  wire nw04548;
  wire nw04549;
  wire nw04550;
  wire nw04551;
  wire nw04552;
  wire nw04553;
  wire nw04554;
  wire nw04555;
  wire nw04556;
  wire nw04557;
  wire nw04558;
  wire nw04559;
  wire nw04560;
  wire nw04561;
  wire nw04562;
  wire nw04563;
  wire nw04564;
  wire nw04565;
  wire nw04566;
  wire nw04567;
  wire nw04568;
  wire nw04569;
  wire nw04570;
  wire nw04571;
  wire nw04572;
  wire nw04573;
  wire nw04574;
  wire nw04575;
  wire nw04576;
  wire nw04577;
  wire nw04578;
  wire nw04579;
  wire nw04580;
  wire nw04581;
  wire nw04582;
  wire nw04583;
  wire nw04584;
  wire nw04585;
  wire nw04586;
  wire nw04587;
  wire nw04588;
  wire nw04589;
  wire nw04590;
  wire nw04591;
  wire nw04592;
  wire nw04593;
  wire nw04594;
  wire nw04595;
  wire nw04596;
  wire nw04597;
  wire nw04598;
  wire nw04599;
  wire nw04600;
  wire nw04601;
  wire nw04602;
  wire nw04603;
  wire nw04604;
  wire nw04605;
  wire nw04606;
  wire nw04607;
  wire nw04608;
  wire nw04609;
  wire nw04610;
  wire nw04611;
  wire nw04612;
  wire nw04613;
  wire nw04614;
  wire nw04615;
  wire nw04616;
  wire nw04617;
  wire nw04618;
  wire nw04619;
  wire nw04620;
  wire nw04621;
  wire nw04622;
  wire nw04623;
  wire nw04624;
  wire nw04625;
  wire nw04626;
  wire nw04627;
  wire nw04628;
  wire nw04629;
  wire nw04630;
  wire nw04631;
  wire nw04632;
  wire nw04633;
  wire nw04634;
  wire nw04635;
  wire nw04636;
  wire nw04637;
  wire nw04638;
  wire nw04639;
  wire nw04640;
  wire nw04641;
  wire nw04642;
  wire nw04643;
  wire nw04644;
  wire nw04645;
  wire nw04646;
  wire nw04647;
  wire nw04648;
  wire nw04649;
  wire nw04650;
  wire nw04651;
  wire nw04652;
  wire nw04653;
  wire nw04654;
  wire nw04655;
  wire nw04656;
  wire nw04657;
  wire nw04658;
  wire nw04659;
  wire nw04660;
  wire nw04661;
  wire nw04662;
  wire nw04663;
  wire nw04664;
  wire nw04665;
  wire nw04666;
  wire nw04667;
  wire nw04668;
  wire nw04669;
  wire nw04670;
  wire nw04671;
  wire nw04672;
  wire nw04673;
  wire nw04674;
  wire nw04675;
  wire nw04676;
  wire nw04677;
  wire nw04678;
  wire nw04679;
  wire nw04680;
  wire nw04681;
  wire nw04682;
  wire nw04683;
  wire nw04684;
  wire nw04685;
  wire nw04686;
  wire nw04687;
  wire nw04688;
  wire nw04689;
  wire nw04690;
  wire nw04691;
  wire nw04692;
  wire nw04693;
  wire nw04694;
  wire nw04695;
  wire nw04696;
  wire nw04697;
  wire nw04698;
  wire nw04699;
  wire nw04700;
  wire nw04701;
  wire nw04702;
  wire nw04703;
  wire nw04704;
  wire nw04705;
  wire nw04706;
  wire nw04707;
  wire nw04708;
  wire nw04709;
  wire nw04710;
  wire nw04711;
  wire nw04712;
  wire nw04713;
  wire nw04714;
  wire nw04715;
  wire nw04716;
  wire nw04717;
  wire nw04718;
  wire nw04719;
  wire nw04720;
  wire nw04721;
  wire nw04722;
  wire nw04723;
  wire nw04724;
  wire nw04725;
  wire nw04726;
  wire nw04727;
  wire nw04728;
  wire nw04729;
  wire nw04730;
  wire nw04731;
  wire nw04732;
  wire nw04733;
  wire nw04734;
  wire nw04735;
  wire nw04736;
  wire nw04737;
  wire nw04738;
  wire nw04739;
  wire nw04740;
  wire nw04741;
  wire nw04742;
  wire nw04743;
  wire nw04744;
  wire nw04745;
  wire nw04746;
  wire nw04747;
  wire nw04748;
  wire nw04749;
  wire nw04750;
  wire nw04751;
  wire nw04752;
  wire nw04753;
  wire nw04754;
  wire nw04755;
  wire nw04756;
  wire nw04757;
  wire nw04758;
  wire nw04759;
  wire nw04760;
  wire nw04761;
  wire nw04762;
  wire nw04763;
  wire nw04764;
  wire nw04765;
  wire nw04766;
  wire nw04767;
  wire nw04768;
  wire nw04769;
  wire nw04770;
  wire nw04771;
  wire nw04772;
  wire nw04773;
  wire nw04774;
  wire nw04775;
  wire nw04776;
  wire nw04777;
  wire nw04778;
  wire nw04779;
  wire nw04780;
  wire nw04781;
  wire nw04782;
  wire nw04783;
  wire nw04784;
  wire nw04785;
  wire nw04786;
  wire nw04787;
  wire nw04788;
  wire nw04789;
  wire nw04790;
  wire nw04791;
  wire nw04792;
  wire nw04793;
  wire nw04794;
  wire nw04795;
  wire nw04796;
  wire nw04797;
  wire nw04798;
  wire nw04799;
  wire nw04800;
  wire nw04801;
  wire nw04802;
  wire nw04803;
  wire nw04804;
  wire nw04805;
  wire nw04806;
  wire nw04807;
  wire nw04808;
  wire nw04809;
  wire nw04810;
  wire nw04811;
  wire nw04812;
  wire nw04813;
  wire nw04814;
  wire nw04815;
  wire nw04816;
  wire nw04817;
  wire nw04818;
  wire nw04819;
  wire nw04820;
  wire nw04821;
  wire nw04822;
  wire nw04823;
  wire nw04824;
  wire nw04825;
  wire nw04826;
  wire nw04827;
  wire nw04828;
  wire nw04829;
  wire nw04830;
  wire nw04831;
  wire nw04832;
  wire nw04833;
  wire nw04834;
  wire nw04835;
  wire nw04836;
  wire nw04837;
  wire nw04838;
  wire nw04839;
  wire nw04840;
  wire nw04841;
  wire nw04842;
  wire nw04843;
  wire nw04844;
  wire nw04845;
  wire nw04846;
  wire nw04847;
  wire nw04848;
  wire nw04849;
  wire nw04850;
  wire nw04851;
  wire nw04852;
  wire nw04853;
  wire nw04854;
  wire nw04855;
  wire nw04856;
  wire nw04857;
  wire nw04858;
  wire nw04859;
  wire nw04860;
  wire nw04861;
  wire nw04862;
  wire nw04863;
  wire nw04864;
  wire nw04865;
  wire nw04866;
  wire nw04867;
  wire nw04868;
  wire nw04869;
  wire nw04870;
  wire nw04871;
  wire nw04872;
  wire nw04873;
  wire nw04874;
  wire nw04875;
  wire nw04876;
  wire nw04877;
  wire nw04878;
  wire nw04879;
  wire nw04880;
  wire nw04881;
  wire nw04882;
  wire nw04883;
  wire nw04884;
  wire nw04885;
  wire nw04886;
  wire nw04887;
  wire nw04888;
  wire nw04889;
  wire nw04890;
  wire nw04891;
  wire nw04892;
  wire nw04893;
  wire nw04894;
  wire nw04895;
  wire nw04896;
  wire nw04897;
  wire nw04898;
  wire nw04899;
  wire nw04900;
  wire nw04901;
  wire nw04902;
  wire nw04903;
  wire nw04904;
  wire nw04905;
  wire nw04906;
  wire nw04907;
  wire nw04908;
  wire nw04909;
  wire nw04910;
  wire nw04911;
  wire nw04912;
  wire nw04913;
  wire nw04914;
  wire nw04915;
  wire nw04916;
  wire nw04917;
  wire nw04918;
  wire nw04919;
  wire nw04920;
  wire nw04921;
  wire nw04922;
  wire nw04923;
  wire nw04924;
  wire nw04925;
  wire nw04926;
  wire nw04927;
  wire nw04928;
  wire nw04929;
  wire nw04930;
  wire nw04931;
  wire nw04932;
  wire nw04933;
  wire nw04934;
  wire nw04935;
  wire nw04936;
  wire nw04937;
  wire nw04938;
  wire nw04939;
  wire nw04940;
  wire nw04941;
  wire nw04942;
  wire nw04943;
  wire nw04944;
  wire nw04945;
  wire nw04946;
  wire nw04947;
  wire nw04948;
  wire nw04949;
  wire nw04950;
  wire nw04951;
  wire nw04952;
  wire nw04953;
  wire nw04954;
  wire nw04955;
  wire nw04956;
  wire nw04957;
  wire nw04958;
  wire nw04959;
  wire nw04960;
  wire nw04961;
  wire nw04962;
  wire nw04963;
  wire nw04964;
  wire nw04965;
  wire nw04966;
  wire nw04967;
  wire nw04968;
  wire nw04969;
  wire nw04970;
  wire nw04971;
  wire nw04972;
  wire nw04973;
  wire nw04974;
  wire nw04975;
  wire nw04976;
  wire nw04977;
  wire nw04978;
  wire nw04979;
  wire nw04980;
  wire nw04981;
  wire nw04982;
  wire nw04983;
  wire nw04984;
  wire nw04985;
  wire nw04986;
  wire nw04987;
  wire nw04988;
  wire nw04989;
  wire nw04990;
  wire nw04991;
  wire nw04992;
  wire nw04993;
  wire nw04994;
  wire nw04995;
  wire nw04996;
  wire nw04997;
  wire nw04998;
  wire nw04999;
  wire nw05000;
  wire nw05001;
  wire nw05002;
  wire nw05003;
  wire nw05004;
  wire nw05005;
  wire nw05006;
  wire nw05007;
  wire nw05008;
  wire nw05009;
  wire nw05010;
  wire nw05011;
  wire nw05012;
  wire nw05013;
  wire nw05014;
  wire nw05015;
  wire nw05016;
  wire nw05017;
  wire nw05018;
  wire nw05019;
  wire nw05020;
  wire nw05021;
  wire nw05022;
  wire nw05023;
  wire nw05024;
  wire nw05025;
  wire nw05026;
  wire nw05027;
  wire nw05028;
  wire nw05029;
  wire nw05030;
  wire nw05031;
  wire nw05032;
  wire nw05033;
  wire nw05034;
  wire nw05035;
  wire nw05036;
  wire nw05037;
  wire nw05038;
  wire nw05039;
  wire nw05040;
  wire nw05041;
  wire nw05042;
  wire nw05043;
  wire nw05044;
  wire nw05045;
  wire nw05046;
  wire nw05047;
  wire nw05048;
  wire nw05049;
  wire nw05050;
  wire nw05051;
  wire nw05052;
  wire nw05053;
  wire nw05054;
  wire nw05055;
  wire nw05056;
  wire nw05057;
  wire nw05058;
  wire nw05059;
  wire nw05060;
  wire nw05061;
  wire nw05062;
  wire nw05063;
  wire nw05064;
  wire nw05065;
  wire nw05066;
  wire nw05067;
  wire nw05068;
  wire nw05069;
  wire nw05070;
  wire nw05071;
  wire nw05072;
  wire nw05073;
  wire nw05074;
  wire nw05075;
  wire nw05076;
  wire nw05077;
  wire nw05078;
  wire nw05079;
  wire nw05080;
  wire nw05081;
  wire nw05082;
  wire nw05083;
  wire nw05084;
  wire nw05085;
  wire nw05086;
  wire nw05087;
  wire nw05088;
  wire nw05089;
  wire nw05090;
  wire nw05091;
  wire nw05092;
  wire nw05093;
  wire nw05094;
  wire nw05095;
  wire nw05096;
  wire nw05097;
  wire nw05098;
  wire nw05099;
  wire nw05100;
  wire nw05101;
  wire nw05102;
  wire nw05103;
  wire nw05104;
  wire nw05105;
  wire nw05106;
  wire nw05107;
  wire nw05108;
  wire nw05109;
  wire nw05110;
  wire nw05111;
  wire nw05112;
  wire nw05113;
  wire nw05114;
  wire nw05115;
  wire nw05116;
  wire nw05117;
  wire nw05118;
  wire nw05119;
  wire nw05120;
  wire nw05121;
  wire nw05122;
  wire nw05123;
  wire nw05124;
  wire nw05125;
  wire nw05126;
  wire nw05127;
  wire nw05128;
  wire nw05129;
  wire nw05130;
  wire nw05131;
  wire nw05132;
  wire nw05133;
  wire nw05134;
  wire nw05135;
  wire nw05136;
  wire nw05137;
  wire nw05138;
  wire nw05139;
  wire nw05140;
  wire nw05141;
  wire nw05142;
  wire nw05143;
  wire nw05144;
  wire nw05145;
  wire nw05146;
  wire nw05147;
  wire nw05148;
  wire nw05149;
  wire nw05150;
  wire nw05151;
  wire nw05152;
  wire nw05153;
  wire nw05154;
  wire nw05155;
  wire nw05156;
  wire nw05157;
  wire nw05158;
  wire nw05159;
  wire nw05160;
  wire nw05161;
  wire nw05162;
  wire nw05163;
  wire nw05164;
  wire nw05165;
  wire nw05166;
  wire nw05167;
  wire nw05168;
  wire nw05169;
  wire nw05170;
  wire nw05171;
  wire nw05172;
  wire nw05173;
  wire nw05174;
  wire nw05175;
  wire nw05176;
  wire nw05177;
  wire nw05178;
  wire nw05179;
  wire nw05180;
  wire nw05181;
  wire nw05182;
  wire nw05183;
  wire nw05184;
  wire nw05185;
  wire nw05186;
  wire nw05187;
  wire nw05188;
  wire nw05189;
  wire nw05190;
  wire nw05191;
  wire nw05192;
  wire nw05193;
  wire nw05194;
  wire nw05195;
  wire nw05196;
  wire nw05197;
  wire nw05198;
  wire nw05199;
  wire nw05200;
  wire nw05201;
  wire nw05202;
  wire nw05203;
  wire nw05204;
  wire nw05205;
  wire nw05206;
  wire nw05207;
  wire nw05208;
  wire nw05209;
  wire nw05210;
  wire nw05211;
  wire nw05212;
  wire nw05213;
  wire nw05214;
  wire nw05215;
  wire nw05216;
  wire nw05217;
  wire nw05218;
  wire nw05219;
  wire nw05220;
  wire nw05221;
  wire nw05222;
  wire nw05223;
  wire nw05224;
  wire nw05225;
  wire nw05226;
  wire nw05227;
  wire nw05228;
  wire nw05229;
  wire nw05230;
  wire nw05231;
  wire nw05232;
  wire nw05233;
  wire nw05234;
  wire nw05235;
  wire nw05236;
  wire nw05237;
  wire nw05238;
  wire nw05239;
  wire nw05240;
  wire nw05241;
  wire nw05242;
  wire nw05243;
  wire nw05244;
  wire nw05245;
  wire nw05246;
  wire nw05247;
  wire nw05248;
  wire nw05249;
  wire nw05250;
  wire nw05251;
  wire nw05252;
  wire nw05253;
  wire nw05254;
  wire nw05255;
  wire nw05256;
  wire nw05257;
  wire nw05258;
  wire nw05259;
  wire nw05260;
  wire nw05261;
  wire nw05262;
  wire nw05263;
  wire nw05264;
  wire nw05265;
  wire nw05266;
  wire nw05267;
  wire nw05268;
  wire nw05269;
  wire nw05270;
  wire nw05271;
  wire nw05272;
  wire nw05273;
  wire nw05274;
  wire nw05275;
  wire nw05276;
  wire nw05277;
  wire nw05278;
  wire nw05279;
  wire nw05280;
  wire nw05281;
  wire nw05282;
  wire nw05283;
  wire nw05284;
  wire nw05285;
  wire nw05286;
  wire nw05287;
  wire nw05288;
  wire nw05289;
  wire nw05290;
  wire nw05291;
  wire nw05292;
  wire nw05293;
  wire nw05294;
  wire nw05295;
  wire nw05296;
  wire nw05297;
  wire nw05298;
  wire nw05299;
  wire nw05300;
  wire nw05301;
  wire nw05302;
  wire nw05303;
  wire nw05304;
  wire nw05305;
  wire nw05306;
  wire nw05307;
  wire nw05308;
  wire nw05309;
  wire nw05310;
  wire nw05311;
  wire nw05312;
  wire nw05313;
  wire nw05314;
  wire nw05315;
  wire nw05316;
  wire nw05317;
  wire nw05318;
  wire nw05319;
  wire nw05320;
  wire nw05321;
  wire nw05322;
  wire nw05323;
  wire nw05324;
  wire nw05325;
  wire nw05326;
  wire nw05327;
  wire nw05328;
  wire nw05329;
  wire nw05330;
  wire nw05331;
  wire nw05332;
  wire nw05333;
  wire nw05334;
  wire nw05335;
  wire nw05336;
  wire nw05337;
  wire nw05338;
  wire nw05339;
  wire nw05340;
  wire nw05341;
  wire nw05342;
  wire nw05343;
  wire nw05344;
  wire nw05345;
  wire nw05346;
  wire nw05347;
  wire nw05348;
  wire nw05349;
  wire nw05350;
  wire nw05351;
  wire nw05352;
  wire nw05353;
  wire nw05354;
  wire nw05355;
  wire nw05356;
  wire nw05357;
  wire nw05358;
  wire nw05359;
  wire nw05360;
  wire nw05361;
  wire nw05362;
  wire nw05363;
  wire nw05364;
  wire nw05365;
  wire nw05366;
  wire nw05367;
  wire nw05368;
  wire nw05369;
  wire nw05370;
  wire nw05371;
  wire nw05372;
  wire nw05373;
  wire nw05374;
  wire nw05375;
  wire nw05376;
  wire nw05377;
  wire nw05378;
  wire nw05379;
  wire nw05380;
  wire nw05381;
  wire nw05382;
  wire nw05383;
  wire nw05384;
  wire nw05385;
  wire nw05386;
  wire nw05387;
  wire nw05388;
  wire nw05389;
  wire nw05390;
  wire nw05391;
  wire nw05392;
  wire nw05393;
  wire nw05394;
  wire nw05395;
  wire nw05396;
  wire nw05397;
  wire nw05398;
  wire nw05399;
  wire nw05400;
  wire nw05401;
  wire nw05402;
  wire nw05403;
  wire nw05404;
  wire nw05405;
  wire nw05406;
  wire nw05407;
  wire nw05408;
  wire [31:0] nw05409;
  wire [31:0] nw05410;
  wire [31:0] nw05411;
  wire [31:0] nw05412;
  wire [31:0] nw05413;
  wire [19:0] nw05414;
  wire [19:0] nw05415;
  wire [3:0] nw05416;
  wire [30:0] nw05417;
  wire [31:0] nw05418;
  wire [31:0] nw05419;
  wire [3:0] nw05420;
  reg [3:0] \nr00002 ;
  reg [3:0] \nr00003 ;
  reg [3:0] \nr00004 ;
  reg [15:0] \nr00005 ;
  reg [15:0] \nr00006 ;
  reg [15:0] \nr00007 ;
  output [31:0] address_ext_o;
  reg [31:0] address_ext_o;
  output [7:0] anodos_o;
  wire [7:0] anodos_o;
  input [3:0] btn_i;
  wire [3:0] btn_i;
  reg nr00008;
  input clock_10_i;
  wire clock_10_i;
  reg [31:0] nr00009;
  wire [31:0] nw05421;
  reg \nr00010 ;
  reg \nr00011 ;
  reg \nr00011u ;
  reg [31:0] \nr00013 ;
  reg [31:0] \nr00014 ;
  reg \nr00015 ;
  reg [31:0] \nr00016 ;
  reg [31:0] \nr00017 ;
  reg [31:0] \nr00018 ;
  reg [31:0] \nr00019 ;
  reg [31:0] \nr00020 ;
  reg [31:0] \nr00021 ;
  reg \nr00021t ;
  reg \nr00021tu ;
  wire [32:0] \nw05422 ;
  reg [31:0] \nr00024 ;
  wire [31:0] \nw05423 ;
  reg [5:0] \nr00025 ;
  wire [31:0] \nw05424 ;
  wire \nw05425 ;
  reg [31:0] \nr00026 ;
  reg \nr00027 ;
  reg \nr00028 ;
  reg \nr00028I ;
  reg \nr00030 ;
  reg \nr00031 ;
  reg \nr00032 ;
  reg \nr00032U ;
  reg \nr00034 ;
  reg \nr00034U ;
  reg \nr00036 ;
  reg \nr00037 ;
  reg \nr00038 ;
  reg \nr00038R ;
  reg \nr00040 ;
  reg \nr00040U ;
  reg \nr00042 ;
  reg \nr00042U ;
  reg \nr00044 ;
  reg \nr00045 ;
  reg \nr00046 ;
  reg \nr00046I ;
  reg \nr00048 ;
  reg \nr00049 ;
  reg \nr00050 ;
  reg \nr00050I ;
  reg \nr00052 ;
  reg \nr00052I ;
  reg \nr00052IU ;
  reg \nr00052U ;
  reg \nr00056 ;
  reg \nr00056I ;
  reg \nr00058 ;
  reg \nr00058I ;
  reg \nr00060 ;
  reg \nr00061 ;
  reg \nr00061I ;
  wire \nw05426 ;
  reg \nr00063 ;
  reg [31:0] \nr00064 ;
  reg \nr00065 ;
  reg [31:0] \nr00066 ;
  reg [31:0] \nr00067 ;
  reg [4:0] \nr00068 ;
  reg [4:0] \nr00069 ;
  reg [4:0] \nr00070 ;
  reg [31:0] \nr00071[0] ;
  reg [31:0] \nr00071[10] ;
  reg [31:0] \nr00071[11] ;
  reg [31:0] \nr00071[12] ;
  reg [31:0] \nr00071[13] ;
  reg [31:0] \nr00071[14] ;
  reg [31:0] \nr00071[15] ;
  reg [31:0] \nr00071[16] ;
  reg [31:0] \nr00071[17] ;
  reg [31:0] \nr00071[18] ;
  reg [31:0] \nr00071[19] ;
  reg [31:0] \nr00071[1] ;
  reg [31:0] \nr00071[20] ;
  reg [31:0] \nr00071[21] ;
  reg [31:0] \nr00071[22] ;
  reg [31:0] \nr00071[23] ;
  reg [31:0] \nr00071[24] ;
  reg [31:0] \nr00071[25] ;
  reg [31:0] \nr00071[26] ;
  reg [31:0] \nr00071[27] ;
  reg [31:0] \nr00071[28] ;
  reg [31:0] \nr00071[29] ;
  reg [31:0] \nr00071[2] ;
  reg [31:0] \nr00071[30] ;
  reg [31:0] \nr00071[31] ;
  reg [31:0] \nr00071[3] ;
  reg [31:0] \nr00071[4] ;
  reg [31:0] \nr00071[5] ;
  reg [31:0] \nr00071[6] ;
  reg [31:0] \nr00071[7] ;
  reg [31:0] \nr00071[8] ;
  reg [31:0] \nr00071[9] ;
  wire [19:0] \nw05427 ;
  reg [3:0] \nr00103  = 4'h0;
  wire \nw05428 ;
  reg [31:0] \nr00104 ;
  output dp_o;
  wire dp_o;
  input [31:0] ext_bus_data_i;
  wire [31:0] ext_bus_data_i;
  output [31:0] ext_bus_data_o;
  reg [31:0] ext_bus_data_o;
  output ext_bus_we_o;
  wire ext_bus_we_o;
  output [10:0] instr_addr_bus_o;
  wire [10:0] instr_addr_bus_o;
  input [31:0] instr_bus_i;
  wire [31:0] instr_bus_i;
  reg [31:0] \nr00105 ;
  wire \nw05429 ;
  output [15:0] led_o;
  wire [15:0] led_o;
  input locked_i;
  wire locked_i;
  output [9:0] ram_address_bus_o;
  wire [9:0] ram_address_bus_o;
  output [31:0] ram_data_in_o;
  wire [31:0] ram_data_in_o;
  input [31:0] ram_data_out_i;
  wire [31:0] ram_data_out_i;
  output ram_we_o;
  wire ram_we_o;
  output reset_effectivo_o;
  wire reset_effectivo_o;
  input reset_i;
  wire reset_i;
  output [6:0] segmentos_o;
  wire [6:0] segmentos_o;
  wire [3:0] nw05430;
  input [15:0] sw_i;
  wire [15:0] sw_i;
  assign nw05414[0] = ~\nw05427 [0];
  assign nw00234 = \nr00016 [0] | \nr00017 [0];
  assign nw05410[0] = \nr00016 [0] & \nr00017 [0];
  assign nw05409[0] = nw00234 & ~(nw05410[0]);
  assign nw00416 = \nr00025 [5] & ~(\nr00063 );
  assign reset_effectivo_o = reset_i | ~(locked_i);
  assign nw00417 = ~(nw05430[2] | nw05430[1]);
  assign nw00418 = ~nw00417;
  assign nw00419 = sw_i[0] | ~(sw_i[1]);
  assign nw00420 = sw_i[3] | sw_i[2];
  assign nw00421 = nw00420 | nw00419;
  assign nw00422 = sw_i[4] | ~(sw_i[5]);
  assign nw00423 = sw_i[7] | sw_i[6];
  assign nw00424 = nw00423 | nw00422;
  assign nw00425 = nw00424 | nw00421;
  assign nw00426 = sw_i[9] | sw_i[8];
  assign nw00427 = sw_i[11] | sw_i[10];
  assign nw00428 = nw00427 | nw00426;
  assign nw00429 = sw_i[12] | ~(sw_i[13]);
  assign nw00430 = sw_i[15] | sw_i[14];
  assign nw00431 = nw00430 | nw00429;
  assign nw00432 = nw00431 | nw00428;
  assign nw00433 = nw00432 | nw00425;
  assign nw00434 = nw05430[0] & ~(nw00433);
  assign nw00435 = nw00434 | nw00418;
  assign nw00436 = ~nw05430[0];
  assign nw00437 = ~(nw00417 & nw00436);
  assign nw00438 = nw00437 & nw00435;
  assign \nw05425  = nw00438 | reset_effectivo_o;
  assign nw00041 = nw00416 & ~(\nw05425 );
  assign nw00439 = ~\nr00063 ;
  assign nw00440 = \nw05425  | nw00439;
  assign nw00441 = \nr00025 [3] & ~(nw00440);
  assign nw00442 = \nw05425  | \nr00063 ;
  assign nw00443 = \nr00025 [0] & ~(nw00442);
  assign nw00003 = nw00443 | nw00441;
  assign nw00444 = ~nw00433;
  assign nw00040 = nw05430[0] ? nw00444 : nw00418;
  assign nw00445 = \nr00025 [2] & ~(nw00440);
  assign nw00446 = \nr00025 [3] & ~(nw00442);
  assign nw00002 = nw00446 | nw00445;
  assign nw00048 = \nr00025 [0] & ~(\nr00063 );
  assign nw00447 = \nr00068 [1] & ~(\nr00068 [0]);
  assign nw00448 = ~(\nr00068 [4] & \nr00068 [3]);
  assign nw00449 = nw00448 | \nr00068 [2];
  assign nw00450 = nw00447 & ~(nw00449);
  assign nw00451 = ~(\nr00025 [4] & \nr00044 );
  assign nw00452 = nw00451 | \nr00063 ;
  assign nw00453 = ~(nw00452 | \nw05425 );
  assign nw00454 = ~\nr00025 [4];
  assign nw00455 = \nr00038R  | \nr00038 ;
  assign nw00456 = \nr00031  | \nr00036 ;
  assign nw00457 = nw00456 | \nr00034 ;
  assign nw00458 = nw00457 | \nr00032 ;
  assign nw00459 = nw00458 | \nr00034U ;
  assign nw00460 = nw00459 | \nr00032U ;
  assign nw00461 = nw00460 | ~(nw00455);
  assign nw00462 = nw00461 | \nr00044 ;
  assign nw00463 = nw00462 | nw00454;
  assign nw00464 = nw00463 | \nr00063 ;
  assign nw00465 = nw00464 | \nw05425 ;
  assign nw00466 = nw00465 & ~(nw00453);
  assign nw00467 = ~\nr00040 ;
  assign nw00468 = address_ext_o[1] | ~(address_ext_o[0]);
  assign nw00469 = nw00468 | nw00467;
  assign nw00470 = nw00469 | nw00455;
  assign nw00471 = nw00470 | nw00460;
  assign nw00472 = nw00471 | \nr00044 ;
  assign nw00473 = nw00472 | nw00454;
  assign nw00474 = nw00473 | \nr00063 ;
  assign nw00475 = ~(nw00474 | \nw05425 );
  assign nw00476 = nw00466 & ~(nw00475);
  assign nw00477 = address_ext_o[0] | ~(address_ext_o[1]);
  assign nw00478 = nw00477 | nw00467;
  assign nw00479 = nw00478 | nw00455;
  assign nw00480 = nw00479 | nw00460;
  assign nw00481 = nw00480 | \nr00044 ;
  assign nw00482 = nw00481 | nw00454;
  assign nw00483 = nw00482 | \nr00063 ;
  assign nw00484 = ~(nw00483 | \nw05425 );
  assign nw00485 = nw00476 & ~(nw00484);
  assign nw00486 = ~(address_ext_o[1] & address_ext_o[0]);
  assign nw00487 = nw00486 | nw00467;
  assign nw00488 = nw00487 | nw00455;
  assign nw00489 = nw00488 | nw00460;
  assign nw00490 = nw00489 | \nr00044 ;
  assign nw00491 = nw00490 | nw00454;
  assign nw00492 = nw00491 | \nr00063 ;
  assign nw00493 = ~(nw00492 | \nw05425 );
  assign nw00494 = nw00485 & ~(nw00493);
  assign nw00495 = address_ext_o[1] | address_ext_o[0];
  assign nw00496 = nw00495 | nw00467;
  assign nw00497 = nw00496 | nw00455;
  assign nw00498 = nw00497 | nw00460;
  assign nw00499 = nw00498 | \nr00044 ;
  assign nw00500 = nw00499 | nw00454;
  assign nw00501 = nw00500 | \nr00063 ;
  assign nw00502 = ~(nw00501 | \nw05425 );
  assign nw00503 = nw00494 & ~(nw00502);
  assign nw00504 = \nr00040  | ~(\nr00042 );
  assign nw00505 = nw00504 | nw00455;
  assign nw00506 = nw00505 | nw00460;
  assign nw00507 = nw00506 | \nr00044 ;
  assign nw00508 = nw00507 | nw00454;
  assign nw00509 = nw00508 | \nr00063 ;
  assign nw00510 = ~(nw00509 | \nw05425 );
  assign nw00511 = nw00503 & ~(nw00510);
  assign nw00512 = \nr00042  | ~(\nr00045 );
  assign nw00513 = nw00512 | \nr00040 ;
  assign nw00514 = nw00513 | nw00455;
  assign nw00515 = nw00514 | nw00460;
  assign nw00516 = nw00515 | \nr00044 ;
  assign nw00517 = nw00516 | nw00454;
  assign nw00518 = nw00517 | \nr00063 ;
  assign nw00519 = ~(nw00518 | \nw05425 );
  assign nw00520 = nw00511 & ~(nw00519);
  assign nw00521 = ~\nr00040U ;
  assign nw00522 = nw00468 | nw00521;
  assign nw00523 = nw00522 | \nr00045 ;
  assign nw00524 = nw00523 | \nr00042 ;
  assign nw00525 = nw00524 | \nr00040 ;
  assign nw00526 = nw00525 | nw00455;
  assign nw00527 = nw00526 | nw00460;
  assign nw00528 = nw00527 | \nr00044 ;
  assign nw00529 = nw00528 | nw00454;
  assign nw00530 = nw00529 | \nr00063 ;
  assign nw00531 = ~(nw00530 | \nw05425 );
  assign nw00532 = nw00520 & ~(nw00531);
  assign nw00533 = nw00477 | nw00521;
  assign nw00534 = nw00533 | \nr00045 ;
  assign nw00535 = nw00534 | \nr00042 ;
  assign nw00536 = nw00535 | \nr00040 ;
  assign nw00537 = nw00536 | nw00455;
  assign nw00538 = nw00537 | nw00460;
  assign nw00539 = nw00538 | \nr00044 ;
  assign nw00540 = nw00539 | nw00454;
  assign nw00541 = nw00540 | \nr00063 ;
  assign nw00542 = ~(nw00541 | \nw05425 );
  assign nw00543 = nw00532 & ~(nw00542);
  assign nw00544 = nw00486 | nw00521;
  assign nw00545 = nw00544 | \nr00045 ;
  assign nw00546 = nw00545 | \nr00042 ;
  assign nw00547 = nw00546 | \nr00040 ;
  assign nw00548 = nw00547 | nw00455;
  assign nw00549 = nw00548 | nw00460;
  assign nw00550 = nw00549 | \nr00044 ;
  assign nw00551 = nw00550 | nw00454;
  assign nw00552 = nw00551 | \nr00063 ;
  assign nw00553 = ~(nw00552 | \nw05425 );
  assign nw00554 = nw00543 & ~(nw00553);
  assign nw00555 = nw00495 | nw00521;
  assign nw00556 = nw00555 | \nr00045 ;
  assign nw00557 = nw00556 | \nr00042 ;
  assign nw00558 = nw00557 | \nr00040 ;
  assign nw00559 = nw00558 | nw00455;
  assign nw00560 = nw00559 | nw00460;
  assign nw00561 = nw00560 | \nr00044 ;
  assign nw00562 = nw00561 | nw00454;
  assign nw00563 = nw00562 | \nr00063 ;
  assign nw00564 = ~(nw00563 | \nw05425 );
  assign nw00565 = nw00554 & ~(nw00564);
  assign nw00566 = \nr00040U  | ~(\nr00042U );
  assign nw00567 = nw00566 | \nr00045 ;
  assign nw00568 = nw00567 | \nr00042 ;
  assign nw00569 = nw00568 | \nr00040 ;
  assign nw00570 = nw00569 | nw00455;
  assign nw00571 = nw00570 | nw00460;
  assign nw00572 = nw00571 | \nr00044 ;
  assign nw00573 = nw00572 | nw00454;
  assign nw00574 = nw00573 | \nr00063 ;
  assign nw00575 = ~(nw00574 | \nw05425 );
  assign nw00576 = nw00565 & ~(nw00575);
  assign nw00577 = \nr00037  | \nr00042U ;
  assign nw00578 = nw00577 | \nr00040U ;
  assign nw00579 = nw00578 | \nr00045 ;
  assign nw00580 = nw00579 | \nr00042 ;
  assign nw00581 = nw00580 | \nr00040 ;
  assign nw00582 = nw00581 | nw00455;
  assign nw00583 = nw00582 | nw00460;
  assign nw00584 = nw00583 | \nr00044 ;
  assign nw00585 = nw00584 | nw00454;
  assign nw00586 = nw00585 | \nr00063 ;
  assign nw00587 = nw00586 | \nw05425 ;
  assign nw00588 = ~(nw00587 & nw00576);
  assign nw00589 = \nr00068 [1] | \nr00068 [0];
  assign nw00590 = \nr00068 [3] | \nr00068 [2];
  assign nw00591 = nw00590 | nw00589;
  assign nw00592 = nw00591 | \nr00068 [4];
  assign nw00593 = ~(nw00592 | \nw05425 );
  assign nw00594 = nw00588 & ~(nw00593);
  assign nw00402 = nw00594 & nw00450;
  assign nw00022 = nw00402 | \nw05425 ;
  assign nw00595 = \nr00010  ? \nr00031  : \nr00036 ;
  assign nw00596 = \nr00034  & ~(\nr00011 );
  assign nw00597 = nw00596 | nw00595;
  assign nw00598 = \nr00032  & \nr00011 ;
  assign nw00599 = nw00598 | nw00597;
  assign nw00600 = \nr00034U  & ~(\nr00011u );
  assign nw00601 = nw00600 | nw00599;
  assign nw00602 = \nr00032U  & \nr00011u ;
  assign nw00603 = nw00602 | nw00601;
  assign nw00604 = \nr00025 [4] & ~(nw00603);
  assign nw00605 = ~\nr00044 ;
  assign nw00606 = ~(nw00460 & nw00605);
  assign nw00607 = nw00604 & ~(nw00606);
  assign nw00608 = nw00451 & ~(nw00607);
  assign nw00609 = \nr00025 [4] & ~(nw00455);
  assign nw00610 = ~nw00609;
  assign nw00611 = nw00460 | nw00467;
  assign nw00612 = nw00611 | nw00610;
  assign nw00613 = nw00605 & ~(nw00612);
  assign nw00614 = nw00460 | ~(\nr00042 );
  assign nw00615 = nw00614 | nw00610;
  assign nw00616 = ~(\nr00044  | \nr00040 );
  assign nw00617 = nw00616 & ~(nw00615);
  assign nw00618 = nw00617 | nw00613;
  assign nw00619 = nw00608 & ~(nw00618);
  assign nw00620 = nw00460 | ~(\nr00045 );
  assign nw00621 = nw00609 & ~(nw00620);
  assign nw00622 = \nr00040  | \nr00042 ;
  assign nw00623 = nw00622 | \nr00044 ;
  assign nw00624 = nw00621 & ~(nw00623);
  assign nw00625 = nw00460 | nw00521;
  assign nw00626 = nw00609 & ~(nw00625);
  assign nw00627 = \nr00042  | \nr00045 ;
  assign nw00628 = nw00627 | ~(nw00616);
  assign nw00629 = nw00626 & ~(nw00628);
  assign nw00630 = nw00629 | nw00624;
  assign nw00631 = nw00460 | ~(\nr00042U );
  assign nw00632 = nw00631 | nw00610;
  assign nw00633 = \nr00045  | \nr00040U ;
  assign nw00634 = nw00633 | nw00622;
  assign nw00635 = nw00634 | nw00632;
  assign nw00636 = nw00605 & ~(nw00635);
  assign nw00637 = nw00460 | \nr00037 ;
  assign nw00638 = nw00637 | nw00610;
  assign nw00639 = \nr00040U  | \nr00042U ;
  assign nw00640 = nw00639 | nw00627;
  assign nw00641 = nw00640 | nw00638;
  assign nw00642 = nw00616 & ~(nw00641);
  assign nw00643 = nw00642 | nw00636;
  assign nw00644 = nw00643 | nw00630;
  assign nw00645 = nw00619 & ~(nw00644);
  assign nw00646 = ~(\nr00025 [0] | \nr00025 [4]);
  assign nw00647 = nw00646 | \nr00063 ;
  assign nw00047 = nw00645 & ~(nw00647);
  assign nw00648 = ~nw00447;
  assign nw00649 = ~\nr00068 [2];
  assign nw00650 = nw00448 | nw00649;
  assign nw00651 = nw00650 | nw00648;
  assign nw00407 = nw00594 & ~(nw00651);
  assign nw00017 = nw00407 | \nw05425 ;
  assign nw00652 = \nr00068 [1] | ~(\nr00068 [0]);
  assign nw00653 = nw00652 | nw00449;
  assign nw00401 = nw00594 & ~(nw00653);
  assign nw00023 = nw00401 | \nw05425 ;
  assign nw00654 = ~(\nr00068 [1] & \nr00068 [0]);
  assign nw00655 = nw00654 | nw00650;
  assign nw00408 = nw00594 & ~(nw00655);
  assign nw00016 = nw00408 | \nw05425 ;
  assign nw00656 = ~(\nr00025 [1] | \nr00025 [0]);
  assign nw00046 = nw00439 & ~(nw00656);
  assign nw00657 = \nr00065  & \nr00063 ;
  assign nw00045 = nw00657 & ~(\nw05425 );
  assign nw00044 = \nr00025 [1] & ~(\nr00063 );
  assign nw00658 = \nr00068 [4] | \nr00068 [3];
  assign nw00659 = nw00658 | \nr00068 [2];
  assign nw00660 = nw00659 | nw00654;
  assign nw00409 = nw00594 & ~(nw00660);
  assign nw00015 = nw00409 | \nw05425 ;
  assign nw00661 = nw00589 | nw00449;
  assign nw00400 = nw00594 & ~(nw00661);
  assign nw00024 = nw00400 | \nw05425 ;
  assign nw00662 = nw00654 | nw00449;
  assign nw00403 = nw00594 & ~(nw00662);
  assign nw00021 = nw00403 | \nw05425 ;
  assign nw00663 = nw00658 | nw00649;
  assign nw00664 = nw00663 | nw00589;
  assign nw00410 = nw00594 & ~(nw00664);
  assign nw00014 = nw00410 | \nw05425 ;
  assign nw00665 = nw00663 | nw00652;
  assign nw00411 = nw00594 & ~(nw00665);
  assign nw00013 = nw00411 | \nw05425 ;
  assign nw00666 = nw00663 | nw00648;
  assign nw00412 = nw00594 & ~(nw00666);
  assign nw00012 = nw00412 | \nw05425 ;
  assign nw00667 = nw00650 | nw00589;
  assign nw00404 = nw00594 & ~(nw00667);
  assign nw00020 = nw00404 | \nw05425 ;
  assign nw00668 = nw00652 | nw00650;
  assign nw00405 = nw00594 & ~(nw00668);
  assign nw00019 = nw00405 | \nw05425 ;
  assign nw00669 = nw00663 | nw00654;
  assign nw00413 = nw00594 & ~(nw00669);
  assign nw00011 = nw00413 | \nw05425 ;
  assign nw00670 = \nr00068 [4] | ~(\nr00068 [3]);
  assign nw00671 = nw00670 | \nr00068 [2];
  assign nw00672 = nw00671 | nw00589;
  assign nw00414 = nw00594 & ~(nw00672);
  assign nw00010 = nw00414 | \nw05425 ;
  assign nw00673 = nw00671 | nw00652;
  assign nw00415 = nw00594 & ~(nw00673);
  assign nw00009 = nw00415 | \nw05425 ;
  assign nw00674 = ~(\nr00013 [0] ^ \nr00014 [0]);
  assign nw00675 = \nr00013 [1] ^ \nr00014 [1];
  assign nw00676 = nw00674 & ~(nw00675);
  assign nw00677 = ~(\nr00013 [3] ^ \nr00014 [3]);
  assign nw00678 = \nr00013 [2] ^ \nr00014 [2];
  assign nw00679 = nw00677 & ~(nw00678);
  assign nw00680 = ~(nw00679 & nw00676);
  assign nw00681 = ~(\nr00013 [7] ^ \nr00014 [7]);
  assign nw00682 = \nr00013 [6] ^ \nr00014 [6];
  assign nw00683 = nw00681 & ~(nw00682);
  assign nw00684 = \nr00013 [5] ^ \nr00014 [5];
  assign nw00685 = \nr00013 [4] ^ \nr00014 [4];
  assign nw00686 = nw00685 | nw00684;
  assign nw00687 = nw00683 & ~(nw00686);
  assign nw00688 = nw00687 & ~(nw00680);
  assign nw00689 = ~(\nr00013 [15] ^ \nr00014 [15]);
  assign nw00690 = \nr00013 [14] ^ \nr00014 [14];
  assign nw00691 = nw00689 & ~(nw00690);
  assign nw00692 = \nr00013 [13] ^ \nr00014 [13];
  assign nw00693 = \nr00013 [12] ^ \nr00014 [12];
  assign nw00694 = nw00693 | nw00692;
  assign nw00695 = nw00691 & ~(nw00694);
  assign nw00696 = ~(\nr00013 [11] ^ \nr00014 [11]);
  assign nw00697 = \nr00013 [10] ^ \nr00014 [10];
  assign nw00698 = nw00696 & ~(nw00697);
  assign nw00699 = \nr00013 [9] ^ \nr00014 [9];
  assign nw00700 = \nr00013 [8] ^ \nr00014 [8];
  assign nw00701 = ~(nw00700 | nw00699);
  assign nw00702 = ~(nw00701 & nw00698);
  assign nw00703 = nw00695 & ~(nw00702);
  assign nw00704 = ~(nw00703 & nw00688);
  assign nw00705 = ~(\nr00013 [31] ^ \nr00014 [31]);
  assign nw00706 = \nr00013 [30] ^ \nr00014 [30];
  assign nw00707 = nw00705 & ~(nw00706);
  assign nw00708 = ~(\nr00013 [29] ^ \nr00014 [29]);
  assign nw00709 = \nr00013 [28] ^ \nr00014 [28];
  assign nw00710 = nw00709 | ~(nw00708);
  assign nw00711 = nw00707 & ~(nw00710);
  assign nw00712 = ~(\nr00013 [27] ^ \nr00014 [27]);
  assign nw00713 = \nr00013 [26] ^ \nr00014 [26];
  assign nw00714 = nw00712 & ~(nw00713);
  assign nw00715 = \nr00013 [25] ^ \nr00014 [25];
  assign nw00716 = \nr00013 [24] ^ \nr00014 [24];
  assign nw00717 = nw00716 | nw00715;
  assign nw00718 = nw00717 | ~(nw00714);
  assign nw00719 = nw00711 & ~(nw00718);
  assign nw00720 = ~(\nr00013 [23] ^ \nr00014 [23]);
  assign nw00721 = \nr00013 [22] ^ \nr00014 [22];
  assign nw00722 = nw00720 & ~(nw00721);
  assign nw00723 = \nr00013 [21] ^ \nr00014 [21];
  assign nw00724 = \nr00013 [20] ^ \nr00014 [20];
  assign nw00725 = nw00724 | nw00723;
  assign nw00726 = nw00722 & ~(nw00725);
  assign nw00727 = ~(\nr00013 [19] ^ \nr00014 [19]);
  assign nw00728 = \nr00013 [18] ^ \nr00014 [18];
  assign nw00729 = nw00727 & ~(nw00728);
  assign nw00730 = \nr00013 [17] ^ \nr00014 [17];
  assign nw00731 = \nr00013 [16] ^ \nr00014 [16];
  assign nw00732 = ~(nw00731 | nw00730);
  assign nw00733 = ~(nw00732 & nw00729);
  assign nw00734 = nw00733 | ~(nw00726);
  assign nw00735 = nw00719 & ~(nw00734);
  assign nw00051 = nw00735 & ~(nw00704);
  assign nw00736 = \nr00013 [31] & ~(\nr00014 [31]);
  assign nw00737 = \nr00014 [30] | ~(\nr00013 [30]);
  assign nw00738 = nw00705 & ~(nw00737);
  assign nw00739 = ~(nw00738 | nw00736);
  assign nw00740 = \nr00014 [29] | ~(\nr00013 [29]);
  assign nw00741 = \nr00014 [28] | ~(\nr00013 [28]);
  assign nw00742 = nw00708 & ~(nw00741);
  assign nw00743 = nw00740 & ~(nw00742);
  assign nw00744 = nw00707 & ~(nw00743);
  assign nw00745 = nw00739 & ~(nw00744);
  assign nw00746 = \nr00014 [27] | ~(\nr00013 [27]);
  assign nw00747 = \nr00014 [26] | ~(\nr00013 [26]);
  assign nw00748 = nw00712 & ~(nw00747);
  assign nw00749 = nw00746 & ~(nw00748);
  assign nw00750 = \nr00014 [25] | ~(\nr00013 [25]);
  assign nw00751 = \nr00013 [24] & ~(\nr00014 [24]);
  assign nw00752 = nw00751 & ~(nw00715);
  assign nw00753 = nw00750 & ~(nw00752);
  assign nw00754 = nw00714 & ~(nw00753);
  assign nw00755 = nw00749 & ~(nw00754);
  assign nw00756 = nw00711 & ~(nw00755);
  assign nw00757 = nw00745 & ~(nw00756);
  assign nw00758 = \nr00014 [23] | ~(\nr00013 [23]);
  assign nw00759 = \nr00014 [22] | ~(\nr00013 [22]);
  assign nw00760 = nw00720 & ~(nw00759);
  assign nw00761 = nw00758 & ~(nw00760);
  assign nw00762 = \nr00014 [21] | ~(\nr00013 [21]);
  assign nw00763 = \nr00013 [20] & ~(\nr00014 [20]);
  assign nw00764 = nw00763 & ~(nw00723);
  assign nw00765 = nw00762 & ~(nw00764);
  assign nw00766 = nw00722 & ~(nw00765);
  assign nw00767 = nw00761 & ~(nw00766);
  assign nw00768 = \nr00014 [19] | ~(\nr00013 [19]);
  assign nw00769 = \nr00014 [18] | ~(\nr00013 [18]);
  assign nw00770 = nw00727 & ~(nw00769);
  assign nw00771 = nw00768 & ~(nw00770);
  assign nw00772 = \nr00014 [17] | ~(\nr00013 [17]);
  assign nw00773 = \nr00013 [16] & ~(\nr00014 [16]);
  assign nw00774 = nw00773 & ~(nw00730);
  assign nw00775 = nw00772 & ~(nw00774);
  assign nw00776 = nw00729 & ~(nw00775);
  assign nw00777 = nw00771 & ~(nw00776);
  assign nw00778 = nw00726 & ~(nw00777);
  assign nw00779 = nw00767 & ~(nw00778);
  assign nw00780 = nw00719 & ~(nw00779);
  assign nw00781 = nw00757 & ~(nw00780);
  assign nw00782 = \nr00014 [15] | ~(\nr00013 [15]);
  assign nw00783 = \nr00014 [14] | ~(\nr00013 [14]);
  assign nw00784 = nw00689 & ~(nw00783);
  assign nw00785 = nw00782 & ~(nw00784);
  assign nw00786 = \nr00014 [13] | ~(\nr00013 [13]);
  assign nw00787 = \nr00013 [12] & ~(\nr00014 [12]);
  assign nw00788 = nw00787 & ~(nw00692);
  assign nw00789 = nw00786 & ~(nw00788);
  assign nw00790 = nw00691 & ~(nw00789);
  assign nw00791 = nw00785 & ~(nw00790);
  assign nw00792 = \nr00014 [11] | ~(\nr00013 [11]);
  assign nw00793 = \nr00014 [10] | ~(\nr00013 [10]);
  assign nw00794 = nw00696 & ~(nw00793);
  assign nw00795 = nw00792 & ~(nw00794);
  assign nw00796 = \nr00014 [9] | ~(\nr00013 [9]);
  assign nw00797 = \nr00013 [8] & ~(\nr00014 [8]);
  assign nw00798 = nw00797 & ~(nw00699);
  assign nw00799 = nw00796 & ~(nw00798);
  assign nw00800 = nw00698 & ~(nw00799);
  assign nw00801 = nw00795 & ~(nw00800);
  assign nw00802 = nw00695 & ~(nw00801);
  assign nw00803 = nw00791 & ~(nw00802);
  assign nw00804 = \nr00014 [7] | ~(\nr00013 [7]);
  assign nw00805 = \nr00014 [6] | ~(\nr00013 [6]);
  assign nw00806 = nw00681 & ~(nw00805);
  assign nw00807 = nw00804 & ~(nw00806);
  assign nw00808 = \nr00014 [5] | ~(\nr00013 [5]);
  assign nw00809 = \nr00013 [4] & ~(\nr00014 [4]);
  assign nw00810 = nw00809 & ~(nw00684);
  assign nw00811 = nw00808 & ~(nw00810);
  assign nw00812 = nw00683 & ~(nw00811);
  assign nw00813 = nw00807 & ~(nw00812);
  assign nw00814 = \nr00014 [3] | ~(\nr00013 [3]);
  assign nw00815 = \nr00014 [2] | ~(\nr00013 [2]);
  assign nw00816 = nw00677 & ~(nw00815);
  assign nw00817 = nw00814 & ~(nw00816);
  assign nw00818 = \nr00014 [1] | ~(\nr00013 [1]);
  assign nw00819 = \nr00013 [0] | ~(\nr00014 [0]);
  assign nw00820 = nw00819 & ~(nw00675);
  assign nw00821 = nw00818 & ~(nw00820);
  assign nw00822 = nw00679 & ~(nw00821);
  assign nw00823 = nw00817 & ~(nw00822);
  assign nw00824 = nw00687 & ~(nw00823);
  assign nw00825 = nw00813 & ~(nw00824);
  assign nw00826 = nw00703 & ~(nw00825);
  assign nw00827 = nw00803 & ~(nw00826);
  assign nw00828 = nw00735 & ~(nw00827);
  assign nw00829 = nw00781 & ~(nw00828);
  assign nw00830 = nw00829 ^ nw00705;
  assign nw00053 = nw00830 | nw00051;
  assign nw00831 = nw00659 | nw00648;
  assign nw00406 = nw00594 & ~(nw00831);
  assign nw00018 = nw00406 | \nw05425 ;
  assign nw00832 = \nr00063  | ~(\nr00025 [3]);
  assign nw00043 = ~(nw00832 | \nw05425 );
  assign nw00052 = nw00051 | ~(nw00829);
  assign nw00833 = \nr00063  | ~(\nr00025 [2]);
  assign nw00042 = ~(nw00833 | \nw05425 );
  assign nw00834 = ~(nr00009[25] | nr00009[24]);
  assign nw00835 = nr00009[27] | nr00009[26];
  assign nw00836 = nw00834 & ~(nw00835);
  assign nw00837 = nr00009[29] | nr00009[28];
  assign nw00838 = nr00009[31] | nr00009[30];
  assign nw00839 = nw00838 | nw00837;
  assign nw00840 = nw00836 & ~(nw00839);
  assign nw00841 = nr00009[23] | nr00009[22];
  assign nw00842 = ~(nr00009[21] | nr00009[20]);
  assign nw00843 = nr00009[23] | ~(nr00009[22]);
  assign nw00844 = nw00842 & ~(nw00843);
  assign nw00845 = nr00009[19] & nr00009[18];
  assign nw00846 = nw00844 & ~(nw00845);
  assign nw00847 = nw00841 & ~(nw00846);
  assign nw00848 = nw00840 & ~(nw00847);
  assign nw00849 = nr00009[17] | nr00009[16];
  assign nw00850 = ~(nr00009[19] & nr00009[18]);
  assign nw00851 = ~(nw00850 | nw00849);
  assign nw00852 = ~(nw00851 & nw00844);
  assign nw00853 = nw00840 & ~(nw00852);
  assign nw00854 = nr00009[15] | nr00009[14];
  assign nw00855 = ~(nr00009[12] | nr00009[13]);
  assign nw00856 = nr00009[15] | ~(nr00009[14]);
  assign nw00857 = nw00855 & ~(nw00856);
  assign nw00858 = nr00009[11] & ~(nr00009[10]);
  assign nw00859 = nr00009[9] & nr00009[8];
  assign nw00860 = nw00858 & ~(nw00859);
  assign nw00861 = nr00009[11] & ~(nw00860);
  assign nw00862 = nw00857 & ~(nw00861);
  assign nw00863 = nw00854 & ~(nw00862);
  assign nw00864 = ~(nr00009[9] & nr00009[8]);
  assign nw00865 = nw00864 | ~(nw00858);
  assign nw00866 = nw00857 & ~(nw00865);
  assign nw00867 = nr00009[7] | nr00009[6];
  assign nw00868 = ~(nr00009[5] | nr00009[4]);
  assign nw00869 = nr00009[7] | ~(nr00009[6]);
  assign nw00870 = nw00868 & ~(nw00869);
  assign nw00871 = nr00009[3] | nr00009[2];
  assign nw00872 = nr00009[1] | nr00009[0];
  assign nw00873 = nw00872 | nw00871;
  assign nw00874 = nw00870 & ~(nw00873);
  assign nw00875 = nw00867 & ~(nw00874);
  assign nw00876 = nw00866 & ~(nw00875);
  assign nw00877 = nw00863 & ~(nw00876);
  assign nw00878 = nw00853 & ~(nw00877);
  assign nw00879 = nw00878 | nw00848;
  assign nw00880 = ~(nw00874 & nw00866);
  assign nw00881 = nw00853 & ~(nw00880);
  assign nw00882 = nw00879 & ~(nw00881);
  assign nw00883 = reset_effectivo_o | ~(nw00882);
  assign nw00884 = nw05430[1] & ~(nw00883);
  assign nw00885 = nw00882 | reset_effectivo_o;
  assign nw00886 = nw05430[2] & ~(nw00885);
  assign nw00007 = nw00886 | nw00884;
  assign nw00887 = nw05430[2] & ~(nw00883);
  assign nw00888 = nw00433 | reset_effectivo_o;
  assign nw00889 = nw00888 | nw00882;
  assign nw00890 = nw05430[0] & ~(nw00889);
  assign nw00008 = nw00890 | nw00887;
  assign nw00891 = \nr00025 [0] & ~(nw00440);
  assign nw00892 = \nr00025 [4] & ~(nw00442);
  assign nw00893 = nw00892 | nw00891;
  assign nw00894 = \nr00048  | \nr00049 ;
  assign nw00895 = ~(nw00894 | \nr00060 );
  assign nw00896 = nw00895 | \nr00063 ;
  assign nw00897 = nw00896 | \nw05425 ;
  assign nw00898 = \nr00025 [1] & ~(nw00897);
  assign nw00899 = nw00898 | \nw05425 ;
  assign nw00000 = nw00899 | nw00893;
  assign nw00900 = nw00888 | ~(nw00882);
  assign nw00901 = nw05430[0] & ~(nw00900);
  assign nw00006 = nw00901 | reset_effectivo_o;
  assign nw00902 = \nr00025 [5] & ~(nw00440);
  assign nw00903 = \nr00025 [2] & ~(nw00442);
  assign nw00005 = nw00903 | nw00902;
  assign nw00904 = \nr00025 [4] & ~(nw00440);
  assign nw00905 = ~(nw00895 & nw00439);
  assign nw00906 = nw00905 | \nw05425 ;
  assign nw00907 = \nr00025 [1] & ~(nw00906);
  assign nw00908 = nw00907 | nw00904;
  assign nw00909 = nw00622 | \nr00045 ;
  assign nw00910 = nw00909 | \nr00040U ;
  assign nw00911 = nw00910 | \nr00042U ;
  assign nw00912 = nw00895 & ~(nw00911);
  assign nw00913 = ~(nw00912 & nw00439);
  assign nw00914 = nw00913 | \nw05425 ;
  assign nw00915 = \nr00025 [5] & ~(nw00914);
  assign nw00004 = nw00915 | nw00908;
  assign nw00916 = \nr00068 [3] | ~(\nr00068 [4]);
  assign nw00917 = nw00916 | nw00649;
  assign nw00918 = nw00917 | nw00652;
  assign nw00397 = nw00594 & ~(nw00918);
  assign nw00027 = nw00397 | \nw05425 ;
  assign nw00919 = nw00917 | nw00648;
  assign nw00398 = nw00594 & ~(nw00919);
  assign nw00026 = nw00398 | \nw05425 ;
  assign nw00920 = nw00917 | nw00654;
  assign nw00399 = nw00594 & ~(nw00920);
  assign nw00025 = nw00399 | \nw05425 ;
  assign nw00921 = \nr00064 [0] & \nr00064 [1];
  assign nw00922 = \nr00064 [3] | ~(\nr00064 [2]);
  assign nw00923 = nw00921 & ~(nw00922);
  assign nw00924 = \nr00064 [5] | ~(\nr00064 [4]);
  assign nw00925 = nw00924 | \nr00064 [6];
  assign nw00103 = nw00923 & ~(nw00925);
  assign nw00926 = ~(\nr00064 [4] & \nr00064 [5]);
  assign nw00927 = nw00926 | \nr00064 [6];
  assign nw00102 = nw00923 & ~(nw00927);
  assign nw00928 = nw00912 | \nr00063 ;
  assign nw00929 = nw00928 | \nw05425 ;
  assign nw00930 = \nr00025 [5] & ~(nw00929);
  assign nw00931 = \nr00025 [1] & ~(nw00440);
  assign nw00001 = nw00931 | nw00930;
  assign nw00932 = nw00917 | nw00589;
  assign nw00396 = nw00594 & ~(nw00932);
  assign nw00028 = nw00396 | \nw05425 ;
  assign nw00933 = nw00659 | nw00652;
  assign nw00395 = nw00594 & ~(nw00933);
  assign nw00029 = nw00395 | \nw05425 ;
  assign nw00934 = nw00916 | \nr00068 [2];
  assign nw00935 = nw00934 | nw00654;
  assign nw00394 = nw00594 & ~(nw00935);
  assign nw00030 = nw00394 | \nw05425 ;
  assign nw00936 = nw00934 | nw00648;
  assign nw00393 = nw00594 & ~(nw00936);
  assign nw00031 = nw00393 | \nw05425 ;
  assign nw00937 = nw00934 | nw00652;
  assign nw00392 = nw00594 & ~(nw00937);
  assign nw00032 = nw00392 | \nw05425 ;
  assign nw00938 = nw00934 | nw00589;
  assign nw00391 = nw00594 & ~(nw00938);
  assign nw00033 = nw00391 | \nw05425 ;
  assign nw00939 = nw00670 | nw00649;
  assign nw00940 = nw00939 | nw00654;
  assign nw00390 = nw00594 & ~(nw00940);
  assign nw00034 = nw00390 | \nw05425 ;
  assign nw00941 = nw00939 | nw00648;
  assign nw00389 = nw00594 & ~(nw00941);
  assign nw00035 = nw00389 | \nw05425 ;
  assign nw00942 = nw00939 | nw00652;
  assign nw00388 = nw00594 & ~(nw00942);
  assign nw00036 = nw00388 | \nw05425 ;
  assign nw00943 = nw00939 | nw00589;
  assign nw00387 = nw00594 & ~(nw00943);
  assign nw00037 = nw00387 | \nw05425 ;
  assign nw00944 = nw00671 | nw00654;
  assign nw00386 = nw00594 & ~(nw00944);
  assign nw00038 = nw00386 | \nw05425 ;
  assign nw00945 = nw00671 | nw00648;
  assign nw00385 = nw00594 & ~(nw00945);
  assign nw00039 = nw00385 | \nw05425 ;
  assign nw00946 = \nr00025 [4] & ~(\nr00044 );
  assign nw00947 = nw00613 | nw00607;
  assign nw00948 = nw00946 & ~(nw00947);
  assign nw00949 = nw00624 | nw00617;
  assign nw00950 = nw00636 | nw00629;
  assign nw00951 = nw00950 | nw00949;
  assign nw00952 = nw00948 & ~(nw00951);
  assign nw00953 = nw00646 | nw00642;
  assign nw00954 = nw00953 | \nr00063 ;
  assign nw00049 = nw00952 & ~(nw00954);
  assign nw00955 = ~(\nr00064 [3] & \nr00064 [2]);
  assign nw00956 = nw00921 & ~(nw00955);
  assign nw00957 = \nr00064 [4] | ~(\nr00064 [5]);
  assign nw00958 = nw00957 | ~(\nr00064 [6]);
  assign nw05416[0] = nw00956 & ~(nw00958);
  assign nw00959 = ~(\nr00064 [3] | \nr00064 [2]);
  assign nw00960 = ~(nw00959 & nw00921);
  assign nw00961 = ~(\nr00064 [12] & \nr00064 [6]);
  assign nw00962 = nw00961 | nw00926;
  assign nw00963 = nw00962 | nw00960;
  assign nw00964 = \nr00064 [14] & ~(\nr00064 [13]);
  assign nw00137 = nw00964 & ~(nw00963);
  assign nw00965 = \nr00064 [12] | \nr00064 [6];
  assign nw00966 = nw00965 | nw00957;
  assign nw00967 = ~(nw00966 | nw00960);
  assign nw00968 = \nr00064 [13] & ~(\nr00064 [14]);
  assign nw00136 = nw00968 & nw00967;
  assign nw00969 = \nr00064 [6] | ~(\nr00064 [12]);
  assign nw00970 = nw00969 | nw00957;
  assign nw00971 = ~(nw00970 | nw00960);
  assign nw00972 = ~(\nr00064 [13] | \nr00064 [14]);
  assign nw00135 = nw00972 & nw00971;
  assign nw00134 = nw00972 & nw00967;
  assign nw00973 = \nr00064 [4] | \nr00064 [5];
  assign nw00974 = nw00973 | nw00969;
  assign nw00975 = nw00974 | nw00960;
  assign nw00133 = nw00964 & ~(nw00975);
  assign nw00976 = nw00973 | nw00965;
  assign nw00977 = nw00976 | nw00960;
  assign nw00132 = nw00964 & ~(nw00977);
  assign nw00131 = nw00968 & ~(nw00977);
  assign nw00130 = nw00972 & ~(nw00975);
  assign nw00129 = nw00972 & ~(nw00977);
  assign nw00978 = ~\nr00064 [31];
  assign nw00979 = nw00969 | nw00926;
  assign nw00980 = nw00979 | nw00960;
  assign nw00981 = \nr00064 [13] & \nr00064 [14];
  assign nw00982 = \nr00064 [26] | \nr00064 [25];
  assign nw00983 = nw00982 | ~(nw00981);
  assign nw00984 = \nr00064 [28] | \nr00064 [27];
  assign nw00985 = \nr00064 [29] | \nr00064 [30];
  assign nw00986 = nw00985 | nw00984;
  assign nw00987 = nw00986 | nw00983;
  assign nw00988 = nw00987 | nw00980;
  assign nw00128 = nw00978 & ~(nw00988);
  assign nw00989 = nw00965 | nw00926;
  assign nw00990 = nw00989 | nw00960;
  assign nw00991 = nw00990 | nw00987;
  assign nw00127 = nw00978 & ~(nw00991);
  assign nw00992 = nw00982 | ~(nw00964);
  assign nw00993 = \nr00064 [29] | ~(\nr00064 [30]);
  assign nw00994 = nw00993 | nw00984;
  assign nw00995 = nw00994 | nw00992;
  assign nw00996 = nw00995 | nw00980;
  assign nw00126 = nw00978 & ~(nw00996);
  assign nw00997 = nw00992 | nw00986;
  assign nw00998 = nw00997 | nw00980;
  assign nw00125 = nw00978 & ~(nw00998);
  assign nw00999 = nw00997 | nw00990;
  assign nw00124 = nw00978 & ~(nw00999);
  assign nw01000 = nw00982 | ~(nw00968);
  assign nw01001 = nw01000 | nw00986;
  assign nw01002 = nw01001 | nw00980;
  assign nw00123 = nw00978 & ~(nw01002);
  assign nw01003 = nw01001 | nw00990;
  assign nw00122 = nw00978 & ~(nw01003);
  assign nw01004 = nw00982 | ~(nw00972);
  assign nw01005 = nw01004 | nw00986;
  assign nw01006 = nw01005 | nw00980;
  assign nw00121 = nw00978 & ~(nw01006);
  assign nw01007 = nw01004 | nw00994;
  assign nw01008 = nw01007 | nw00990;
  assign nw00120 = nw00978 & ~(nw01008);
  assign nw01009 = nw01005 | nw00990;
  assign nw00119 = nw00978 & ~(nw01009);
  assign nw01010 = nw00969 | nw00924;
  assign nw01011 = nw01010 | nw00960;
  assign nw01012 = nw01011 | nw00995;
  assign nw00118 = nw00978 & ~(nw01012);
  assign nw01013 = nw01011 | nw00997;
  assign nw00117 = nw00978 & ~(nw01013);
  assign nw01014 = nw01011 | nw01005;
  assign nw00116 = nw00978 & ~(nw01014);
  assign nw00115 = nw00981 & ~(nw01011);
  assign nw01015 = nw00965 | nw00924;
  assign nw01016 = nw01015 | nw00960;
  assign nw00114 = nw00981 & ~(nw01016);
  assign nw00113 = nw00964 & ~(nw01016);
  assign nw00112 = nw00968 & ~(nw01011);
  assign nw00111 = nw00968 & ~(nw01016);
  assign nw01017 = nw00961 | nw00957;
  assign nw01018 = nw01017 | nw00960;
  assign nw00110 = nw00981 & ~(nw01018);
  assign nw01019 = \nr00064 [12] | ~(\nr00064 [6]);
  assign nw01020 = nw01019 | nw00957;
  assign nw01021 = nw01020 | nw00960;
  assign nw00109 = nw00981 & ~(nw01021);
  assign nw00108 = nw00964 & ~(nw01018);
  assign nw00107 = nw00964 & ~(nw01021);
  assign nw00106 = nw00972 & ~(nw01018);
  assign nw00105 = nw00972 & ~(nw01021);
  assign nw01022 = nw01020 | ~(nw00923);
  assign nw00104 = nw00972 & ~(nw01022);
  assign nw05421[0] = nw00882 & ~(nr00009[0]);
  assign nw01023 = ~(nr00009[1] ^ nr00009[0]);
  assign nw05421[1] = nw00882 & ~(nw01023);
  assign nw01024 = nr00009[1] & nr00009[0];
  assign nw01025 = ~(nw01024 ^ nr00009[2]);
  assign nw05421[2] = nw00882 & ~(nw01025);
  assign nw01026 = ~(nw01024 & nr00009[2]);
  assign nw01027 = nw01026 ^ nr00009[3];
  assign nw05421[3] = nw00882 & ~(nw01027);
  assign nw01028 = ~(nr00009[3] & nr00009[2]);
  assign nw01029 = nw01024 & ~(nw01028);
  assign nw01030 = ~(nw01029 ^ nr00009[4]);
  assign nw05421[4] = nw00882 & ~(nw01030);
  assign nw01031 = ~(nw01029 & nr00009[4]);
  assign nw01032 = nw01031 ^ nr00009[5];
  assign nw05421[5] = nw00882 & ~(nw01032);
  assign nw01033 = ~(nr00009[5] & nr00009[4]);
  assign nw01034 = nw01029 & ~(nw01033);
  assign nw01035 = ~(nw01034 ^ nr00009[6]);
  assign nw05421[6] = nw00882 & ~(nw01035);
  assign nw01036 = ~(nw01034 & nr00009[6]);
  assign nw01037 = nw01036 ^ nr00009[7];
  assign nw05421[7] = nw00882 & ~(nw01037);
  assign nw01038 = ~(nr00009[7] & nr00009[6]);
  assign nw01039 = ~(nw01038 | nw01033);
  assign nw01040 = ~(nw01039 & nw01029);
  assign nw01041 = nw01040 ^ nr00009[8];
  assign nw05421[8] = nw00882 & ~(nw01041);
  assign nw01042 = nw01040 | ~(nr00009[8]);
  assign nw01043 = nw01042 ^ nr00009[9];
  assign nw05421[9] = nw00882 & ~(nw01043);
  assign nw01044 = ~(nw01040 | nw00864);
  assign nw01045 = ~(nw01044 ^ nr00009[10]);
  assign nw05421[10] = nw00882 & ~(nw01045);
  assign nw01046 = ~(nw01044 & nr00009[10]);
  assign nw01047 = nw01046 ^ nr00009[11];
  assign nw05421[11] = nw00882 & ~(nw01047);
  assign nw01048 = ~(nr00009[10] & nr00009[11]);
  assign nw01049 = nw01048 | nw00864;
  assign nw01050 = ~(nw01049 | nw01040);
  assign nw01051 = ~(nw01050 ^ nr00009[12]);
  assign nw05421[12] = nw00882 & ~(nw01051);
  assign nw01052 = ~(nw01050 & nr00009[12]);
  assign nw01053 = nw01052 ^ nr00009[13];
  assign nw05421[13] = nw00882 & ~(nw01053);
  assign nw01054 = ~(nr00009[12] & nr00009[13]);
  assign nw01055 = nw01050 & ~(nw01054);
  assign nw01056 = ~(nw01055 ^ nr00009[14]);
  assign nw05421[14] = nw00882 & ~(nw01056);
  assign nw01057 = ~(nw01055 & nr00009[14]);
  assign nw01058 = nw01057 ^ nr00009[15];
  assign nw05421[15] = nw00882 & ~(nw01058);
  assign nw01059 = ~(nr00009[15] & nr00009[14]);
  assign nw01060 = nw01059 | nw01054;
  assign nw01061 = nw01060 | nw01049;
  assign nw01062 = ~(nw01061 | nw01040);
  assign nw01063 = ~(nw01062 ^ nr00009[16]);
  assign nw05421[16] = nw00882 & ~(nw01063);
  assign nw01064 = ~(nw01062 & nr00009[16]);
  assign nw01065 = nw01064 ^ nr00009[17];
  assign nw05421[17] = nw00882 & ~(nw01065);
  assign nw01066 = ~(nr00009[17] & nr00009[16]);
  assign nw01067 = nw01062 & ~(nw01066);
  assign nw01068 = ~(nw01067 ^ nr00009[18]);
  assign nw05421[18] = nw00882 & ~(nw01068);
  assign nw01069 = ~(nw01067 & nr00009[18]);
  assign nw01070 = nw01069 ^ nr00009[19];
  assign nw05421[19] = nw00882 & ~(nw01070);
  assign nw01071 = nw01066 | nw00850;
  assign nw01072 = nw01062 & ~(nw01071);
  assign nw01073 = ~(nw01072 ^ nr00009[20]);
  assign nw05421[20] = nw00882 & ~(nw01073);
  assign nw01074 = ~(nw01072 & nr00009[20]);
  assign nw01075 = nw01074 ^ nr00009[21];
  assign nw05421[21] = nw00882 & ~(nw01075);
  assign nw01076 = ~(nr00009[21] & nr00009[20]);
  assign nw01077 = nw01072 & ~(nw01076);
  assign nw01078 = ~(nw01077 ^ nr00009[22]);
  assign nw05421[22] = nw00882 & ~(nw01078);
  assign nw01079 = ~(nw01077 & nr00009[22]);
  assign nw01080 = nw01079 ^ nr00009[23];
  assign nw05421[23] = nw00882 & ~(nw01080);
  assign nw01081 = ~(nr00009[23] & nr00009[22]);
  assign nw01082 = nw01081 | nw01076;
  assign nw01083 = nw01082 | nw01071;
  assign nw01084 = nw01062 & ~(nw01083);
  assign nw01085 = ~(nw01084 ^ nr00009[24]);
  assign nw05421[24] = nw00882 & ~(nw01085);
  assign nw01086 = ~(nw01084 & nr00009[24]);
  assign nw01087 = nw01086 ^ nr00009[25];
  assign nw05421[25] = nw00882 & ~(nw01087);
  assign nw01088 = ~(nr00009[25] & nr00009[24]);
  assign nw01089 = nw01084 & ~(nw01088);
  assign nw01090 = ~(nw01089 ^ nr00009[26]);
  assign nw05421[26] = nw00882 & ~(nw01090);
  assign nw01091 = ~(nw01089 & nr00009[26]);
  assign nw01092 = nw01091 ^ nr00009[27];
  assign nw05421[27] = nw00882 & ~(nw01092);
  assign nw01093 = ~(nr00009[27] & nr00009[26]);
  assign nw01094 = nw01093 | nw01088;
  assign nw01095 = nw01084 & ~(nw01094);
  assign nw01096 = ~(nw01095 ^ nr00009[28]);
  assign nw05421[28] = nw00882 & ~(nw01096);
  assign nw01097 = ~(nw01095 & nr00009[28]);
  assign nw01098 = nw01097 ^ nr00009[29];
  assign nw05421[29] = nw00882 & ~(nw01098);
  assign nw01099 = ~(nr00009[29] & nr00009[28]);
  assign nw01100 = nw01095 & ~(nw01099);
  assign nw01101 = ~(nw01100 ^ nr00009[30]);
  assign nw05421[30] = nw00882 & ~(nw01101);
  assign nw01102 = ~(nw01100 & nr00009[30]);
  assign nw01103 = nw01102 ^ nr00009[31];
  assign nw05421[31] = nw00882 & ~(nw01103);
  assign nw01104 = address_ext_o[31] | address_ext_o[30];
  assign nw01105 = address_ext_o[29] | address_ext_o[28];
  assign nw01106 = nw01105 | nw01104;
  assign nw01107 = address_ext_o[27] | address_ext_o[26];
  assign nw01108 = address_ext_o[25] | address_ext_o[24];
  assign nw01109 = nw01108 | nw01107;
  assign nw01110 = nw01109 | nw01106;
  assign nw01111 = address_ext_o[23] | address_ext_o[22];
  assign nw01112 = address_ext_o[21] | address_ext_o[20];
  assign nw01113 = nw01112 | nw01111;
  assign nw01114 = address_ext_o[19] | address_ext_o[18];
  assign nw01115 = address_ext_o[17] | address_ext_o[16];
  assign nw01116 = nw01115 | nw01114;
  assign nw01117 = nw01116 | nw01113;
  assign nw01118 = nw01117 | nw01110;
  assign nw01119 = ~(address_ext_o[15] | address_ext_o[14]);
  assign nw01120 = ~(address_ext_o[13] | address_ext_o[12]);
  assign nw01121 = ~(nw01120 & nw01119);
  assign nw01122 = nw01121 | address_ext_o[11];
  assign nw01123 = address_ext_o[7] | address_ext_o[6];
  assign nw01124 = address_ext_o[5] | address_ext_o[4];
  assign nw01125 = nw01124 | nw01123;
  assign nw01126 = address_ext_o[2] | address_ext_o[3];
  assign nw01127 = nw00495 | nw01126;
  assign nw01128 = nw01127 | nw01125;
  assign nw01129 = address_ext_o[9] | address_ext_o[8];
  assign nw01130 = address_ext_o[10] | ~(address_ext_o[11]);
  assign nw01131 = nw01130 | nw01129;
  assign nw01132 = nw01131 | nw01121;
  assign nw01133 = ~(nw01132 | nw01128);
  assign nw01134 = nw01122 & ~(nw01133);
  assign nw01135 = ~(nw01134 | nw01118);
  assign nw01136 = nw01133 & ~(nw01118);
  assign nw01137 = nw01135 & ~(nw01136);
  assign nw01138 = ~(address_ext_o[11] | address_ext_o[10]);
  assign nw01139 = nw01129 | ~(nw01138);
  assign nw01140 = address_ext_o[13] & ~(address_ext_o[12]);
  assign nw01141 = ~(nw01140 & nw01119);
  assign nw01142 = nw01141 | nw01139;
  assign nw01143 = address_ext_o[3] | ~(address_ext_o[2]);
  assign nw01144 = nw01143 | nw00495;
  assign nw01145 = nw01144 | nw01125;
  assign nw01146 = nw01145 | nw01142;
  assign nw01147 = ~(nw01146 | nw01118);
  assign nw01148 = address_ext_o[2] | ~(address_ext_o[3]);
  assign nw01149 = nw01148 | nw00495;
  assign nw01150 = nw01149 | nw01125;
  assign nw01151 = nw01150 | nw01142;
  assign nw01152 = ~(nw01151 | nw01118);
  assign nw01153 = address_ext_o[5] | ~(address_ext_o[4]);
  assign nw01154 = nw01153 | nw01123;
  assign nw01155 = nw01154 | nw01127;
  assign nw01156 = nw01155 | nw01142;
  assign nw01157 = ~(nw01156 | nw01118);
  assign nw01158 = address_ext_o[13] & address_ext_o[12];
  assign nw01159 = ~(nw01158 & nw01119);
  assign nw01160 = nw01159 | nw01139;
  assign nw01161 = nw01160 | nw01128;
  assign nw01162 = nw01161 | nw01118;
  assign nw01163 = nw01119 & ~(nw01158);
  assign nw01164 = nw01161 & ~(nw01163);
  assign nw01165 = nw01164 | nw01118;
  assign nw01166 = nw01162 & ~(nw01165);
  assign nw01167 = nw01160 & ~(nw01163);
  assign nw01168 = address_ext_o[8] & ~(address_ext_o[9]);
  assign nw01169 = ~(nw01168 & nw01138);
  assign nw01170 = nw01169 | nw01159;
  assign nw01171 = ~(nw01170 | nw01128);
  assign nw01172 = nw01167 & ~(nw01171);
  assign nw01173 = nw01172 | nw01118;
  assign nw01174 = nw01171 & ~(nw01118);
  assign nw01175 = nw01174 | nw01173;
  assign nw01176 = nw01175 | nw01166;
  assign nw01177 = ext_bus_data_i[0] & ~(nw01176);
  assign nw01178 = nw01157 ? \nr00007 [0] : nw01177;
  assign nw01179 = nw01152 ? \nr00104 [0] : nw01178;
  assign nw01180 = nw01147 ? \nr00105 [0] : nw01179;
  assign nw01181 = address_ext_o[12] & ~(address_ext_o[13]);
  assign nw01182 = ~(nw01181 & nw01119);
  assign nw01183 = nw01182 | nw01139;
  assign nw01184 = nw01183 | nw01128;
  assign nw01185 = ~(nw01184 | nw01118);
  assign nw01186 = nw01184 & nw01121;
  assign nw01187 = nw01186 | nw01118;
  assign nw01188 = nw01187 | nw01185;
  assign nw01189 = nw01138 & ~(nw01182);
  assign nw01190 = nw01121 & ~(nw01189);
  assign nw01191 = address_ext_o[11] | ~(address_ext_o[10]);
  assign nw01192 = nw01191 | nw01129;
  assign nw01193 = nw01192 | nw01182;
  assign nw01194 = ~(nw01193 | nw01128);
  assign nw01195 = nw01190 & ~(nw01194);
  assign nw01196 = nw01195 | nw01118;
  assign nw01197 = nw01194 & ~(nw01118);
  assign nw01198 = nw01197 | nw01196;
  assign nw01199 = nw01188 & ~(nw01198);
  assign nw01200 = nw01199 ? ram_data_out_i[0] : nw01180;
  assign \nw05424 [0] = nw01137 ? instr_bus_i[0] : nw01200;
  assign nw01201 = ext_bus_data_i[1] & ~(nw01176);
  assign nw01202 = nw01157 ? \nr00007 [1] : nw01201;
  assign nw01203 = nw01152 ? \nr00104 [1] : nw01202;
  assign nw01204 = nw01147 ? \nr00105 [1] : nw01203;
  assign nw01205 = nw01199 ? ram_data_out_i[1] : nw01204;
  assign \nw05424 [1] = nw01137 ? instr_bus_i[1] : nw01205;
  assign nw01206 = ext_bus_data_i[2] & ~(nw01176);
  assign nw01207 = nw01157 ? \nr00007 [2] : nw01206;
  assign nw01208 = nw01152 ? \nr00104 [2] : nw01207;
  assign nw01209 = nw01147 ? \nr00105 [2] : nw01208;
  assign nw01210 = nw01199 ? ram_data_out_i[2] : nw01209;
  assign \nw05424 [2] = nw01137 ? instr_bus_i[2] : nw01210;
  assign nw01211 = ext_bus_data_i[3] & ~(nw01176);
  assign nw01212 = nw01157 ? \nr00007 [3] : nw01211;
  assign nw01213 = nw01152 ? \nr00104 [3] : nw01212;
  assign nw01214 = nw01147 ? \nr00105 [3] : nw01213;
  assign nw01215 = nw01199 ? ram_data_out_i[3] : nw01214;
  assign \nw05424 [3] = nw01137 ? instr_bus_i[3] : nw01215;
  assign nw01216 = ext_bus_data_i[4] & ~(nw01176);
  assign nw01217 = nw01157 ? \nr00007 [4] : nw01216;
  assign nw01218 = nw01152 ? \nr00104 [4] : nw01217;
  assign nw01219 = nw01147 ? \nr00105 [4] : nw01218;
  assign nw01220 = nw01199 ? ram_data_out_i[4] : nw01219;
  assign \nw05424 [4] = nw01137 ? instr_bus_i[4] : nw01220;
  assign nw01221 = ext_bus_data_i[5] & ~(nw01176);
  assign nw01222 = nw01157 ? \nr00007 [5] : nw01221;
  assign nw01223 = nw01152 ? \nr00104 [5] : nw01222;
  assign nw01224 = nw01147 ? \nr00105 [5] : nw01223;
  assign nw01225 = nw01199 ? ram_data_out_i[5] : nw01224;
  assign \nw05424 [5] = nw01137 ? instr_bus_i[5] : nw01225;
  assign nw01226 = ext_bus_data_i[6] & ~(nw01176);
  assign nw01227 = nw01157 ? \nr00007 [6] : nw01226;
  assign nw01228 = nw01152 ? \nr00104 [6] : nw01227;
  assign nw01229 = nw01147 ? \nr00105 [6] : nw01228;
  assign nw01230 = nw01199 ? ram_data_out_i[6] : nw01229;
  assign \nw05424 [6] = nw01137 ? instr_bus_i[6] : nw01230;
  assign nw01231 = ext_bus_data_i[7] & ~(nw01176);
  assign nw01232 = nw01157 ? \nr00007 [7] : nw01231;
  assign nw01233 = nw01152 ? \nr00104 [7] : nw01232;
  assign nw01234 = nw01147 ? \nr00105 [7] : nw01233;
  assign nw01235 = nw01199 ? ram_data_out_i[7] : nw01234;
  assign \nw05424 [7] = nw01137 ? instr_bus_i[7] : nw01235;
  assign nw01236 = ext_bus_data_i[8] & ~(nw01176);
  assign nw01237 = nw01157 ? \nr00007 [8] : nw01236;
  assign nw01238 = nw01152 ? \nr00104 [8] : nw01237;
  assign nw01239 = nw01147 ? \nr00105 [8] : nw01238;
  assign nw01240 = nw01199 ? ram_data_out_i[8] : nw01239;
  assign \nw05424 [8] = nw01137 ? instr_bus_i[8] : nw01240;
  assign nw01241 = ext_bus_data_i[9] & ~(nw01176);
  assign nw01242 = nw01157 ? \nr00007 [9] : nw01241;
  assign nw01243 = nw01152 ? \nr00104 [9] : nw01242;
  assign nw01244 = nw01147 ? \nr00105 [9] : nw01243;
  assign nw01245 = nw01199 ? ram_data_out_i[9] : nw01244;
  assign \nw05424 [9] = nw01137 ? instr_bus_i[9] : nw01245;
  assign nw01246 = ext_bus_data_i[10] & ~(nw01176);
  assign nw01247 = nw01157 ? \nr00007 [10] : nw01246;
  assign nw01248 = nw01152 ? \nr00104 [10] : nw01247;
  assign nw01249 = nw01147 ? \nr00105 [10] : nw01248;
  assign nw01250 = nw01199 ? ram_data_out_i[10] : nw01249;
  assign \nw05424 [10] = nw01137 ? instr_bus_i[10] : nw01250;
  assign nw01251 = ext_bus_data_i[11] & ~(nw01176);
  assign nw01252 = nw01157 ? \nr00007 [11] : nw01251;
  assign nw01253 = nw01152 ? \nr00104 [11] : nw01252;
  assign nw01254 = nw01147 ? \nr00105 [11] : nw01253;
  assign nw01255 = nw01199 ? ram_data_out_i[11] : nw01254;
  assign \nw05424 [11] = nw01137 ? instr_bus_i[11] : nw01255;
  assign nw01256 = ext_bus_data_i[12] & ~(nw01176);
  assign nw01257 = nw01157 ? \nr00007 [12] : nw01256;
  assign nw01258 = nw01152 ? \nr00104 [12] : nw01257;
  assign nw01259 = nw01147 ? \nr00105 [12] : nw01258;
  assign nw01260 = nw01199 ? ram_data_out_i[12] : nw01259;
  assign \nw05424 [12] = nw01137 ? instr_bus_i[12] : nw01260;
  assign nw01261 = ext_bus_data_i[13] & ~(nw01176);
  assign nw01262 = nw01157 ? \nr00007 [13] : nw01261;
  assign nw01263 = nw01152 ? \nr00104 [13] : nw01262;
  assign nw01264 = nw01147 ? \nr00105 [13] : nw01263;
  assign nw01265 = nw01199 ? ram_data_out_i[13] : nw01264;
  assign \nw05424 [13] = nw01137 ? instr_bus_i[13] : nw01265;
  assign nw01266 = ext_bus_data_i[14] & ~(nw01176);
  assign nw01267 = nw01157 ? \nr00007 [14] : nw01266;
  assign nw01268 = nw01152 ? \nr00104 [14] : nw01267;
  assign nw01269 = nw01147 ? \nr00105 [14] : nw01268;
  assign nw01270 = nw01199 ? ram_data_out_i[14] : nw01269;
  assign \nw05424 [14] = nw01137 ? instr_bus_i[14] : nw01270;
  assign nw01271 = ext_bus_data_i[15] & ~(nw01176);
  assign nw01272 = nw01157 ? \nr00007 [15] : nw01271;
  assign nw01273 = nw01152 ? \nr00104 [15] : nw01272;
  assign nw01274 = nw01147 ? \nr00105 [15] : nw01273;
  assign nw01275 = nw01199 ? ram_data_out_i[15] : nw01274;
  assign \nw05424 [15] = nw01137 ? instr_bus_i[15] : nw01275;
  assign nw01276 = ext_bus_data_i[16] & ~(nw01176);
  assign nw01277 = nw01157 ? \nr00004 [0] : nw01276;
  assign nw01278 = nw01152 ? \nr00104 [16] : nw01277;
  assign nw01279 = nw01147 ? \nr00105 [16] : nw01278;
  assign nw01280 = nw01199 ? ram_data_out_i[16] : nw01279;
  assign \nw05424 [16] = nw01137 ? instr_bus_i[16] : nw01280;
  assign nw01281 = ext_bus_data_i[17] & ~(nw01176);
  assign nw01282 = nw01157 ? \nr00004 [1] : nw01281;
  assign nw01283 = nw01152 ? \nr00104 [17] : nw01282;
  assign nw01284 = nw01147 ? \nr00105 [17] : nw01283;
  assign nw01285 = nw01199 ? ram_data_out_i[17] : nw01284;
  assign \nw05424 [17] = nw01137 ? instr_bus_i[17] : nw01285;
  assign nw01286 = ext_bus_data_i[18] & ~(nw01176);
  assign nw01287 = nw01157 ? \nr00004 [2] : nw01286;
  assign nw01288 = nw01152 ? \nr00104 [18] : nw01287;
  assign nw01289 = nw01147 ? \nr00105 [18] : nw01288;
  assign nw01290 = nw01199 ? ram_data_out_i[18] : nw01289;
  assign \nw05424 [18] = nw01137 ? instr_bus_i[18] : nw01290;
  assign nw01291 = ext_bus_data_i[19] & ~(nw01176);
  assign nw01292 = nw01157 ? \nr00004 [3] : nw01291;
  assign nw01293 = nw01152 ? \nr00104 [19] : nw01292;
  assign nw01294 = nw01147 ? \nr00105 [19] : nw01293;
  assign nw01295 = nw01199 ? ram_data_out_i[19] : nw01294;
  assign \nw05424 [19] = nw01137 ? instr_bus_i[19] : nw01295;
  assign nw01296 = nw01176 | ~(ext_bus_data_i[20]);
  assign nw01297 = ~(nw01296 | nw01157);
  assign nw01298 = nw01152 ? \nr00104 [20] : nw01297;
  assign nw01299 = nw01147 ? \nr00105 [20] : nw01298;
  assign nw01300 = nw01199 ? ram_data_out_i[20] : nw01299;
  assign \nw05424 [20] = nw01137 ? instr_bus_i[20] : nw01300;
  assign nw01301 = nw01176 | ~(ext_bus_data_i[21]);
  assign nw01302 = ~(nw01301 | nw01157);
  assign nw01303 = nw01152 ? \nr00104 [21] : nw01302;
  assign nw01304 = nw01147 ? \nr00105 [21] : nw01303;
  assign nw01305 = nw01199 ? ram_data_out_i[21] : nw01304;
  assign \nw05424 [21] = nw01137 ? instr_bus_i[21] : nw01305;
  assign nw01306 = nw01176 | ~(ext_bus_data_i[22]);
  assign nw01307 = ~(nw01306 | nw01157);
  assign nw01308 = nw01152 ? \nr00104 [22] : nw01307;
  assign nw01309 = nw01147 ? \nr00105 [22] : nw01308;
  assign nw01310 = nw01199 ? ram_data_out_i[22] : nw01309;
  assign \nw05424 [22] = nw01137 ? instr_bus_i[22] : nw01310;
  assign nw01311 = nw01176 | ~(ext_bus_data_i[23]);
  assign nw01312 = ~(nw01311 | nw01157);
  assign nw01313 = nw01152 ? \nr00104 [23] : nw01312;
  assign nw01314 = nw01147 ? \nr00105 [23] : nw01313;
  assign nw01315 = nw01199 ? ram_data_out_i[23] : nw01314;
  assign \nw05424 [23] = nw01137 ? instr_bus_i[23] : nw01315;
  assign nw01316 = nw01176 | ~(ext_bus_data_i[24]);
  assign nw01317 = ~(nw01316 | nw01157);
  assign nw01318 = nw01152 ? \nr00104 [24] : nw01317;
  assign nw01319 = nw01147 ? \nr00105 [24] : nw01318;
  assign nw01320 = nw01199 ? ram_data_out_i[24] : nw01319;
  assign \nw05424 [24] = nw01137 ? instr_bus_i[24] : nw01320;
  assign nw01321 = nw01176 | ~(ext_bus_data_i[25]);
  assign nw01322 = ~(nw01321 | nw01157);
  assign nw01323 = nw01152 ? \nr00104 [25] : nw01322;
  assign nw01324 = nw01147 ? \nr00105 [25] : nw01323;
  assign nw01325 = nw01199 ? ram_data_out_i[25] : nw01324;
  assign \nw05424 [25] = nw01137 ? instr_bus_i[25] : nw01325;
  assign nw01326 = nw01176 | ~(ext_bus_data_i[26]);
  assign nw01327 = ~(nw01326 | nw01157);
  assign nw01328 = nw01152 ? \nr00104 [26] : nw01327;
  assign nw01329 = nw01147 ? \nr00105 [26] : nw01328;
  assign nw01330 = nw01199 ? ram_data_out_i[26] : nw01329;
  assign \nw05424 [26] = nw01137 ? instr_bus_i[26] : nw01330;
  assign nw01331 = nw01176 | ~(ext_bus_data_i[27]);
  assign nw01332 = ~(nw01331 | nw01157);
  assign nw01333 = nw01152 ? \nr00104 [27] : nw01332;
  assign nw01334 = nw01147 ? \nr00105 [27] : nw01333;
  assign nw01335 = nw01199 ? ram_data_out_i[27] : nw01334;
  assign \nw05424 [27] = nw01137 ? instr_bus_i[27] : nw01335;
  assign nw01336 = nw01176 | ~(ext_bus_data_i[28]);
  assign nw01337 = ~(nw01336 | nw01157);
  assign nw01338 = nw01152 ? \nr00104 [28] : nw01337;
  assign nw01339 = nw01147 ? \nr00105 [28] : nw01338;
  assign nw01340 = nw01199 ? ram_data_out_i[28] : nw01339;
  assign \nw05424 [28] = nw01137 ? instr_bus_i[28] : nw01340;
  assign nw01341 = nw01176 | ~(ext_bus_data_i[29]);
  assign nw01342 = ~(nw01341 | nw01157);
  assign nw01343 = nw01152 ? \nr00104 [29] : nw01342;
  assign nw01344 = nw01147 ? \nr00105 [29] : nw01343;
  assign nw01345 = nw01199 ? ram_data_out_i[29] : nw01344;
  assign \nw05424 [29] = nw01137 ? instr_bus_i[29] : nw01345;
  assign nw01346 = nw01176 | ~(ext_bus_data_i[30]);
  assign nw01347 = ~(nw01346 | nw01157);
  assign nw01348 = nw01152 ? \nr00104 [30] : nw01347;
  assign nw01349 = nw01147 ? \nr00105 [30] : nw01348;
  assign nw01350 = nw01199 ? ram_data_out_i[30] : nw01349;
  assign \nw05424 [30] = nw01137 ? instr_bus_i[30] : nw01350;
  assign nw01351 = nw01176 | ~(ext_bus_data_i[31]);
  assign nw01352 = ~(nw01351 | nw01157);
  assign nw01353 = nw01152 ? \nr00104 [31] : nw01352;
  assign nw01354 = nw01147 ? \nr00105 [31] : nw01353;
  assign nw01355 = nw01199 ? ram_data_out_i[31] : nw01354;
  assign \nw05424 [31] = nw01137 ? instr_bus_i[31] : nw01355;
  assign nw01356 = ~(nw01152 & nr00008);
  assign nw01357 = nw01356 | nw01147;
  assign \nw05428  = ~(nw01357 | nw01199);
  assign nw01358 = ~(nw01147 & nr00008);
  assign \nw05429  = ~(nw01358 | nw01199);
  assign nw01359 = address_ext_o[1] ? \nr00064 [16] : \nr00064 [0];
  assign nw01360 = nw00465 ? \nr00026 [0] : \nr00066 [0];
  assign nw01361 = nw00475 ? \nr00064 [8] : nw01360;
  assign nw01362 = nw00484 ? \nr00064 [16] : nw01361;
  assign nw01363 = nw00493 ? \nr00064 [24] : nw01362;
  assign nw01364 = nw00502 ? \nr00064 [0] : nw01363;
  assign nw01365 = nw00510 ? nw01359 : nw01364;
  assign nw01366 = nw00519 ? \nr00064 [0] : nw01365;
  assign nw01367 = nw00531 ? \nr00064 [8] : nw01366;
  assign nw01368 = nw00542 ? \nr00064 [16] : nw01367;
  assign nw01369 = nw00553 ? \nr00064 [24] : nw01368;
  assign nw01370 = nw00564 ? \nr00064 [0] : nw01369;
  assign nw01371 = nw00575 ? nw01359 : nw01370;
  assign nw01372 = \nr00015  ? \nr00024 [0] : \nr00018 [0];
  assign nw01373 = ~(\nr00056I  | \nr00056 );
  assign nw01374 = \nr00058  | ~(nw01373);
  assign nw01375 = nw01374 | \nr00058I ;
  assign nw01376 = nw01375 ? \nw05422 [0] : nw01372;
  assign nw01377 = \nr00050I  | \nr00050 ;
  assign nw01378 = nw01377 ? \nr00021 [0] : nw01376;
  assign nw01379 = \nr00028I  | \nr00028 ;
  assign nw01380 = nw01379 ? \nr00019 [0] : nw01378;
  assign nw01381 = \nr00046I  | \nr00046 ;
  assign nw01382 = nw01381 ? \nr00020 [0] : nw01380;
  assign nw01383 = \nr00061I  | \nr00061 ;
  assign nw01384 = nw01383 ? \nr00018 [0] : nw01382;
  assign nw01385 = \nr00052IU  | \nr00052U ;
  assign nw01386 = nw01385 ? \nr00021tu  : nw01384;
  assign nw01387 = \nr00052I  | \nr00052 ;
  assign nw01388 = nw01387 ? \nr00021t  : nw01386;
  assign nw00065 = nw00587 ? nw01371 : nw01388;
  assign nw01389 = address_ext_o[1] ? \nr00064 [17] : \nr00064 [1];
  assign nw01390 = nw00465 ? \nr00026 [1] : \nr00066 [1];
  assign nw01391 = nw00475 ? \nr00064 [9] : nw01390;
  assign nw01392 = nw00484 ? \nr00064 [17] : nw01391;
  assign nw01393 = nw00493 ? \nr00064 [25] : nw01392;
  assign nw01394 = nw00502 ? \nr00064 [1] : nw01393;
  assign nw01395 = nw00510 ? nw01389 : nw01394;
  assign nw01396 = nw00519 ? \nr00064 [1] : nw01395;
  assign nw01397 = nw00531 ? \nr00064 [9] : nw01396;
  assign nw01398 = nw00542 ? \nr00064 [17] : nw01397;
  assign nw01399 = nw00553 ? \nr00064 [25] : nw01398;
  assign nw01400 = nw00564 ? \nr00064 [1] : nw01399;
  assign nw01401 = nw00575 ? nw01389 : nw01400;
  assign nw01402 = ~\nw05423 [1];
  assign nw01403 = ~\nr00020 [1];
  assign nw01404 = ~\nr00019 [1];
  assign nw01405 = ~\nr00021 [1];
  assign nw01406 = ~\nw05422 [1];
  assign nw01407 = ~\nr00018 [1];
  assign nw01408 = ~\nr00024 [1];
  assign nw01409 = \nr00015  ? nw01408 : nw01407;
  assign nw01410 = nw01375 ? nw01406 : nw01409;
  assign nw01411 = nw01377 ? nw01405 : nw01410;
  assign nw01412 = nw01379 ? nw01404 : nw01411;
  assign nw01413 = nw01381 ? nw01403 : nw01412;
  assign nw01414 = nw01383 ? nw01402 : nw01413;
  assign nw01415 = nw01414 | nw01385;
  assign nw01416 = ~(nw01415 | nw01387);
  assign nw00076 = nw00587 ? nw01401 : nw01416;
  assign nw01417 = address_ext_o[1] ? \nr00064 [18] : \nr00064 [2];
  assign nw01418 = nw00465 ? \nr00026 [2] : \nr00066 [2];
  assign nw01419 = nw00475 ? \nr00064 [10] : nw01418;
  assign nw01420 = nw00484 ? \nr00064 [18] : nw01419;
  assign nw01421 = nw00493 ? \nr00064 [26] : nw01420;
  assign nw01422 = nw00502 ? \nr00064 [2] : nw01421;
  assign nw01423 = nw00510 ? nw01417 : nw01422;
  assign nw01424 = nw00519 ? \nr00064 [2] : nw01423;
  assign nw01425 = nw00531 ? \nr00064 [10] : nw01424;
  assign nw01426 = nw00542 ? \nr00064 [18] : nw01425;
  assign nw01427 = nw00553 ? \nr00064 [26] : nw01426;
  assign nw01428 = nw00564 ? \nr00064 [2] : nw01427;
  assign nw01429 = nw00575 ? nw01417 : nw01428;
  assign nw01430 = ~\nw05423 [2];
  assign nw01431 = ~\nr00020 [2];
  assign nw01432 = ~\nr00019 [2];
  assign nw01433 = ~\nr00021 [2];
  assign nw01434 = ~\nw05422 [2];
  assign nw01435 = ~\nr00018 [2];
  assign nw01436 = ~\nr00024 [2];
  assign nw01437 = \nr00015  ? nw01436 : nw01435;
  assign nw01438 = nw01375 ? nw01434 : nw01437;
  assign nw01439 = nw01377 ? nw01433 : nw01438;
  assign nw01440 = nw01379 ? nw01432 : nw01439;
  assign nw01441 = nw01381 ? nw01431 : nw01440;
  assign nw01442 = nw01383 ? nw01430 : nw01441;
  assign nw01443 = nw01442 | nw01385;
  assign nw01444 = ~(nw01443 | nw01387);
  assign nw00087 = nw00587 ? nw01429 : nw01444;
  assign nw01445 = address_ext_o[1] ? \nr00064 [19] : \nr00064 [3];
  assign nw01446 = nw00465 ? \nr00026 [3] : \nr00066 [3];
  assign nw01447 = nw00475 ? \nr00064 [11] : nw01446;
  assign nw01448 = nw00484 ? \nr00064 [19] : nw01447;
  assign nw01449 = nw00493 ? \nr00064 [27] : nw01448;
  assign nw01450 = nw00502 ? \nr00064 [3] : nw01449;
  assign nw01451 = nw00510 ? nw01445 : nw01450;
  assign nw01452 = nw00519 ? \nr00064 [3] : nw01451;
  assign nw01453 = nw00531 ? \nr00064 [11] : nw01452;
  assign nw01454 = nw00542 ? \nr00064 [19] : nw01453;
  assign nw01455 = nw00553 ? \nr00064 [27] : nw01454;
  assign nw01456 = nw00564 ? \nr00064 [3] : nw01455;
  assign nw01457 = nw00575 ? nw01445 : nw01456;
  assign nw01458 = ~\nw05423 [3];
  assign nw01459 = ~\nr00020 [3];
  assign nw01460 = ~\nr00019 [3];
  assign nw01461 = ~\nr00021 [3];
  assign nw01462 = ~\nw05422 [3];
  assign nw01463 = ~\nr00018 [3];
  assign nw01464 = ~\nr00024 [3];
  assign nw01465 = \nr00015  ? nw01464 : nw01463;
  assign nw01466 = nw01375 ? nw01462 : nw01465;
  assign nw01467 = nw01377 ? nw01461 : nw01466;
  assign nw01468 = nw01379 ? nw01460 : nw01467;
  assign nw01469 = nw01381 ? nw01459 : nw01468;
  assign nw01470 = nw01383 ? nw01458 : nw01469;
  assign nw01471 = nw01470 | nw01385;
  assign nw01472 = ~(nw01471 | nw01387);
  assign nw00090 = nw00587 ? nw01457 : nw01472;
  assign nw01473 = address_ext_o[1] ? \nr00064 [20] : \nr00064 [4];
  assign nw01474 = nw00465 ? \nr00026 [4] : \nr00066 [4];
  assign nw01475 = nw00475 ? \nr00064 [12] : nw01474;
  assign nw01476 = nw00484 ? \nr00064 [20] : nw01475;
  assign nw01477 = nw00493 ? \nr00064 [28] : nw01476;
  assign nw01478 = nw00502 ? \nr00064 [4] : nw01477;
  assign nw01479 = nw00510 ? nw01473 : nw01478;
  assign nw01480 = nw00519 ? \nr00064 [4] : nw01479;
  assign nw01481 = nw00531 ? \nr00064 [12] : nw01480;
  assign nw01482 = nw00542 ? \nr00064 [20] : nw01481;
  assign nw01483 = nw00553 ? \nr00064 [28] : nw01482;
  assign nw01484 = nw00564 ? \nr00064 [4] : nw01483;
  assign nw01485 = nw00575 ? nw01473 : nw01484;
  assign nw01486 = ~\nw05423 [4];
  assign nw01487 = ~\nr00020 [4];
  assign nw01488 = ~\nr00019 [4];
  assign nw01489 = ~\nr00021 [4];
  assign nw01490 = ~\nw05422 [4];
  assign nw01491 = ~\nr00018 [4];
  assign nw01492 = ~\nr00024 [4];
  assign nw01493 = \nr00015  ? nw01492 : nw01491;
  assign nw01494 = nw01375 ? nw01490 : nw01493;
  assign nw01495 = nw01377 ? nw01489 : nw01494;
  assign nw01496 = nw01379 ? nw01488 : nw01495;
  assign nw01497 = nw01381 ? nw01487 : nw01496;
  assign nw01498 = nw01383 ? nw01486 : nw01497;
  assign nw01499 = nw01498 | nw01385;
  assign nw01500 = ~(nw01499 | nw01387);
  assign nw00091 = nw00587 ? nw01485 : nw01500;
  assign nw01501 = address_ext_o[1] ? \nr00064 [21] : \nr00064 [5];
  assign nw01502 = nw00465 ? \nr00026 [5] : \nr00066 [5];
  assign nw01503 = nw00475 ? \nr00064 [13] : nw01502;
  assign nw01504 = nw00484 ? \nr00064 [21] : nw01503;
  assign nw01505 = nw00493 ? \nr00064 [29] : nw01504;
  assign nw01506 = nw00502 ? \nr00064 [5] : nw01505;
  assign nw01507 = nw00510 ? nw01501 : nw01506;
  assign nw01508 = nw00519 ? \nr00064 [5] : nw01507;
  assign nw01509 = nw00531 ? \nr00064 [13] : nw01508;
  assign nw01510 = nw00542 ? \nr00064 [21] : nw01509;
  assign nw01511 = nw00553 ? \nr00064 [29] : nw01510;
  assign nw01512 = nw00564 ? \nr00064 [5] : nw01511;
  assign nw01513 = nw00575 ? nw01501 : nw01512;
  assign nw01514 = ~\nw05423 [5];
  assign nw01515 = ~\nr00020 [5];
  assign nw01516 = ~\nr00019 [5];
  assign nw01517 = ~\nr00021 [5];
  assign nw01518 = ~\nw05422 [5];
  assign nw01519 = ~\nr00018 [5];
  assign nw01520 = ~\nr00024 [5];
  assign nw01521 = \nr00015  ? nw01520 : nw01519;
  assign nw01522 = nw01375 ? nw01518 : nw01521;
  assign nw01523 = nw01377 ? nw01517 : nw01522;
  assign nw01524 = nw01379 ? nw01516 : nw01523;
  assign nw01525 = nw01381 ? nw01515 : nw01524;
  assign nw01526 = nw01383 ? nw01514 : nw01525;
  assign nw01527 = nw01526 | nw01385;
  assign nw01528 = ~(nw01527 | nw01387);
  assign nw00092 = nw00587 ? nw01513 : nw01528;
  assign nw01529 = address_ext_o[1] ? \nr00064 [22] : \nr00064 [6];
  assign nw01530 = nw00465 ? \nr00026 [6] : \nr00066 [6];
  assign nw01531 = nw00475 ? \nr00064 [14] : nw01530;
  assign nw01532 = nw00484 ? \nr00064 [22] : nw01531;
  assign nw01533 = nw00493 ? \nr00064 [30] : nw01532;
  assign nw01534 = nw00502 ? \nr00064 [6] : nw01533;
  assign nw01535 = nw00510 ? nw01529 : nw01534;
  assign nw01536 = nw00519 ? \nr00064 [6] : nw01535;
  assign nw01537 = nw00531 ? \nr00064 [14] : nw01536;
  assign nw01538 = nw00542 ? \nr00064 [22] : nw01537;
  assign nw01539 = nw00553 ? \nr00064 [30] : nw01538;
  assign nw01540 = nw00564 ? \nr00064 [6] : nw01539;
  assign nw01541 = nw00575 ? nw01529 : nw01540;
  assign nw01542 = ~\nw05423 [6];
  assign nw01543 = ~\nr00020 [6];
  assign nw01544 = ~\nr00019 [6];
  assign nw01545 = ~\nr00021 [6];
  assign nw01546 = ~\nw05422 [6];
  assign nw01547 = ~\nr00018 [6];
  assign nw01548 = ~\nr00024 [6];
  assign nw01549 = \nr00015  ? nw01548 : nw01547;
  assign nw01550 = nw01375 ? nw01546 : nw01549;
  assign nw01551 = nw01377 ? nw01545 : nw01550;
  assign nw01552 = nw01379 ? nw01544 : nw01551;
  assign nw01553 = nw01381 ? nw01543 : nw01552;
  assign nw01554 = nw01383 ? nw01542 : nw01553;
  assign nw01555 = nw01554 | nw01385;
  assign nw01556 = ~(nw01555 | nw01387);
  assign nw00093 = nw00587 ? nw01541 : nw01556;
  assign nw01557 = address_ext_o[1] ? \nr00064 [23] : \nr00064 [7];
  assign nw01558 = nw00465 ? \nr00026 [7] : \nr00066 [7];
  assign nw01559 = nw00475 ? \nr00064 [15] : nw01558;
  assign nw01560 = nw00484 ? \nr00064 [23] : nw01559;
  assign nw01561 = nw00493 ? \nr00064 [31] : nw01560;
  assign nw01562 = nw00502 ? \nr00064 [7] : nw01561;
  assign nw01563 = nw00510 ? nw01557 : nw01562;
  assign nw01564 = nw00519 ? \nr00064 [7] : nw01563;
  assign nw01565 = nw00531 ? \nr00064 [15] : nw01564;
  assign nw01566 = nw00542 ? \nr00064 [23] : nw01565;
  assign nw01567 = nw00553 ? \nr00064 [31] : nw01566;
  assign nw01568 = nw00564 ? \nr00064 [7] : nw01567;
  assign nw01569 = nw00575 ? nw01557 : nw01568;
  assign nw01570 = ~\nw05423 [7];
  assign nw01571 = ~\nr00020 [7];
  assign nw01572 = ~\nr00019 [7];
  assign nw01573 = ~\nr00021 [7];
  assign nw01574 = ~\nw05422 [7];
  assign nw01575 = ~\nr00018 [7];
  assign nw01576 = ~\nr00024 [7];
  assign nw01577 = \nr00015  ? nw01576 : nw01575;
  assign nw01578 = nw01375 ? nw01574 : nw01577;
  assign nw01579 = nw01377 ? nw01573 : nw01578;
  assign nw01580 = nw01379 ? nw01572 : nw01579;
  assign nw01581 = nw01381 ? nw01571 : nw01580;
  assign nw01582 = nw01383 ? nw01570 : nw01581;
  assign nw01583 = nw01582 | nw01385;
  assign nw01584 = ~(nw01583 | nw01387);
  assign nw00094 = nw00587 ? nw01569 : nw01584;
  assign nw01585 = ~\nr00064 [8];
  assign nw01586 = ~\nr00064 [24];
  assign nw01587 = address_ext_o[1] ? nw01586 : nw01585;
  assign nw01588 = ~nw01587;
  assign nw01589 = ~\nr00064 [7];
  assign nw01590 = ~\nr00064 [23];
  assign nw01591 = ~\nr00064 [15];
  assign nw01592 = ~\nr00026 [8];
  assign nw01593 = ~\nr00066 [8];
  assign nw01594 = nw00465 ? nw01592 : nw01593;
  assign nw01595 = nw00475 ? nw01591 : nw01594;
  assign nw01596 = nw00484 ? nw01590 : nw01595;
  assign nw01597 = nw00493 ? nw00978 : nw01596;
  assign nw01598 = nw00502 ? nw01589 : nw01597;
  assign nw01599 = nw00510 ? nw01587 : nw01598;
  assign nw01600 = nw00519 ? nw01585 : nw01599;
  assign nw01601 = nw01600 | nw00531;
  assign nw01602 = nw01601 | nw00542;
  assign nw01603 = nw01602 | nw00553;
  assign nw01604 = ~(nw01603 | nw00564);
  assign nw01605 = nw00575 ? nw01588 : nw01604;
  assign nw01606 = ~\nw05423 [8];
  assign nw01607 = ~\nr00020 [8];
  assign nw01608 = ~\nr00019 [8];
  assign nw01609 = ~\nr00021 [8];
  assign nw01610 = ~\nw05422 [8];
  assign nw01611 = ~\nr00018 [8];
  assign nw01612 = ~\nr00024 [8];
  assign nw01613 = \nr00015  ? nw01612 : nw01611;
  assign nw01614 = nw01375 ? nw01610 : nw01613;
  assign nw01615 = nw01377 ? nw01609 : nw01614;
  assign nw01616 = nw01379 ? nw01608 : nw01615;
  assign nw01617 = nw01381 ? nw01607 : nw01616;
  assign nw01618 = nw01383 ? nw01606 : nw01617;
  assign nw01619 = nw01618 | nw01385;
  assign nw01620 = ~(nw01619 | nw01387);
  assign nw00095 = nw00587 ? nw01605 : nw01620;
  assign nw01621 = ~\nr00064 [25];
  assign nw01622 = ~\nr00064 [9];
  assign nw01623 = address_ext_o[1] ? nw01621 : nw01622;
  assign nw01624 = ~nw01623;
  assign nw01625 = ~\nr00026 [9];
  assign nw01626 = ~\nr00066 [9];
  assign nw01627 = nw00465 ? nw01625 : nw01626;
  assign nw01628 = nw00475 ? nw01591 : nw01627;
  assign nw01629 = nw00484 ? nw01590 : nw01628;
  assign nw01630 = nw00493 ? nw00978 : nw01629;
  assign nw01631 = nw00502 ? nw01589 : nw01630;
  assign nw01632 = nw00510 ? nw01623 : nw01631;
  assign nw01633 = nw00519 ? nw01622 : nw01632;
  assign nw01634 = nw01633 | nw00531;
  assign nw01635 = nw01634 | nw00542;
  assign nw01636 = nw01635 | nw00553;
  assign nw01637 = ~(nw01636 | nw00564);
  assign nw01638 = nw00575 ? nw01624 : nw01637;
  assign nw01639 = ~\nw05423 [9];
  assign nw01640 = ~\nr00020 [9];
  assign nw01641 = ~\nr00019 [9];
  assign nw01642 = ~\nr00021 [9];
  assign nw01643 = ~\nw05422 [9];
  assign nw01644 = ~\nr00018 [9];
  assign nw01645 = ~\nr00024 [9];
  assign nw01646 = \nr00015  ? nw01645 : nw01644;
  assign nw01647 = nw01375 ? nw01643 : nw01646;
  assign nw01648 = nw01377 ? nw01642 : nw01647;
  assign nw01649 = nw01379 ? nw01641 : nw01648;
  assign nw01650 = nw01381 ? nw01640 : nw01649;
  assign nw01651 = nw01383 ? nw01639 : nw01650;
  assign nw01652 = nw01651 | nw01385;
  assign nw01653 = ~(nw01652 | nw01387);
  assign nw00096 = nw00587 ? nw01638 : nw01653;
  assign nw01654 = ~\nr00064 [26];
  assign nw01655 = ~\nr00064 [10];
  assign nw01656 = address_ext_o[1] ? nw01654 : nw01655;
  assign nw01657 = ~nw01656;
  assign nw01658 = ~\nr00026 [10];
  assign nw01659 = ~\nr00066 [10];
  assign nw01660 = nw00465 ? nw01658 : nw01659;
  assign nw01661 = nw00475 ? nw01591 : nw01660;
  assign nw01662 = nw00484 ? nw01590 : nw01661;
  assign nw01663 = nw00493 ? nw00978 : nw01662;
  assign nw01664 = nw00502 ? nw01589 : nw01663;
  assign nw01665 = nw00510 ? nw01656 : nw01664;
  assign nw01666 = nw00519 ? nw01655 : nw01665;
  assign nw01667 = nw01666 | nw00531;
  assign nw01668 = nw01667 | nw00542;
  assign nw01669 = nw01668 | nw00553;
  assign nw01670 = ~(nw01669 | nw00564);
  assign nw01671 = nw00575 ? nw01657 : nw01670;
  assign nw01672 = ~\nw05423 [10];
  assign nw01673 = ~\nr00020 [10];
  assign nw01674 = ~\nr00019 [10];
  assign nw01675 = ~\nr00021 [10];
  assign nw01676 = ~\nw05422 [10];
  assign nw01677 = ~\nr00018 [10];
  assign nw01678 = ~\nr00024 [10];
  assign nw01679 = \nr00015  ? nw01678 : nw01677;
  assign nw01680 = nw01375 ? nw01676 : nw01679;
  assign nw01681 = nw01377 ? nw01675 : nw01680;
  assign nw01682 = nw01379 ? nw01674 : nw01681;
  assign nw01683 = nw01381 ? nw01673 : nw01682;
  assign nw01684 = nw01383 ? nw01672 : nw01683;
  assign nw01685 = nw01684 | nw01385;
  assign nw01686 = ~(nw01685 | nw01387);
  assign nw00066 = nw00587 ? nw01671 : nw01686;
  assign nw01687 = ~\nr00064 [27];
  assign nw01688 = ~\nr00064 [11];
  assign nw01689 = address_ext_o[1] ? nw01687 : nw01688;
  assign nw01690 = ~nw01689;
  assign nw01691 = ~\nr00026 [11];
  assign nw01692 = ~\nr00066 [11];
  assign nw01693 = nw00465 ? nw01691 : nw01692;
  assign nw01694 = nw00475 ? nw01591 : nw01693;
  assign nw01695 = nw00484 ? nw01590 : nw01694;
  assign nw01696 = nw00493 ? nw00978 : nw01695;
  assign nw01697 = nw00502 ? nw01589 : nw01696;
  assign nw01698 = nw00510 ? nw01689 : nw01697;
  assign nw01699 = nw00519 ? nw01688 : nw01698;
  assign nw01700 = nw01699 | nw00531;
  assign nw01701 = nw01700 | nw00542;
  assign nw01702 = nw01701 | nw00553;
  assign nw01703 = ~(nw01702 | nw00564);
  assign nw01704 = nw00575 ? nw01690 : nw01703;
  assign nw01705 = ~\nw05423 [11];
  assign nw01706 = ~\nr00020 [11];
  assign nw01707 = ~\nr00019 [11];
  assign nw01708 = ~\nr00021 [11];
  assign nw01709 = ~\nw05422 [11];
  assign nw01710 = ~\nr00018 [11];
  assign nw01711 = ~\nr00024 [11];
  assign nw01712 = \nr00015  ? nw01711 : nw01710;
  assign nw01713 = nw01375 ? nw01709 : nw01712;
  assign nw01714 = nw01377 ? nw01708 : nw01713;
  assign nw01715 = nw01379 ? nw01707 : nw01714;
  assign nw01716 = nw01381 ? nw01706 : nw01715;
  assign nw01717 = nw01383 ? nw01705 : nw01716;
  assign nw01718 = nw01717 | nw01385;
  assign nw01719 = ~(nw01718 | nw01387);
  assign nw00067 = nw00587 ? nw01704 : nw01719;
  assign nw01720 = ~\nr00064 [12];
  assign nw01721 = ~\nr00064 [28];
  assign nw01722 = address_ext_o[1] ? nw01721 : nw01720;
  assign nw01723 = ~nw01722;
  assign nw01724 = ~\nr00026 [12];
  assign nw01725 = ~\nr00066 [12];
  assign nw01726 = nw00465 ? nw01724 : nw01725;
  assign nw01727 = nw00475 ? nw01591 : nw01726;
  assign nw01728 = nw00484 ? nw01590 : nw01727;
  assign nw01729 = nw00493 ? nw00978 : nw01728;
  assign nw01730 = nw00502 ? nw01589 : nw01729;
  assign nw01731 = nw00510 ? nw01722 : nw01730;
  assign nw01732 = nw00519 ? nw01720 : nw01731;
  assign nw01733 = nw01732 | nw00531;
  assign nw01734 = nw01733 | nw00542;
  assign nw01735 = nw01734 | nw00553;
  assign nw01736 = ~(nw01735 | nw00564);
  assign nw01737 = nw00575 ? nw01723 : nw01736;
  assign nw01738 = ~\nw05423 [12];
  assign nw01739 = ~\nr00020 [12];
  assign nw01740 = ~\nr00019 [12];
  assign nw01741 = ~\nr00021 [12];
  assign nw01742 = ~\nw05422 [12];
  assign nw01743 = ~\nr00018 [12];
  assign nw01744 = ~\nr00024 [12];
  assign nw01745 = \nr00015  ? nw01744 : nw01743;
  assign nw01746 = nw01375 ? nw01742 : nw01745;
  assign nw01747 = nw01377 ? nw01741 : nw01746;
  assign nw01748 = nw01379 ? nw01740 : nw01747;
  assign nw01749 = nw01381 ? nw01739 : nw01748;
  assign nw01750 = nw01383 ? nw01738 : nw01749;
  assign nw01751 = nw01750 | nw01385;
  assign nw01752 = ~(nw01751 | nw01387);
  assign nw00068 = nw00587 ? nw01737 : nw01752;
  assign nw01753 = ~\nr00064 [13];
  assign nw01754 = ~\nr00064 [29];
  assign nw01755 = address_ext_o[1] ? nw01754 : nw01753;
  assign nw01756 = ~nw01755;
  assign nw01757 = ~\nr00026 [13];
  assign nw01758 = ~\nr00066 [13];
  assign nw01759 = nw00465 ? nw01757 : nw01758;
  assign nw01760 = nw00475 ? nw01591 : nw01759;
  assign nw01761 = nw00484 ? nw01590 : nw01760;
  assign nw01762 = nw00493 ? nw00978 : nw01761;
  assign nw01763 = nw00502 ? nw01589 : nw01762;
  assign nw01764 = nw00510 ? nw01755 : nw01763;
  assign nw01765 = nw00519 ? nw01753 : nw01764;
  assign nw01766 = nw01765 | nw00531;
  assign nw01767 = nw01766 | nw00542;
  assign nw01768 = nw01767 | nw00553;
  assign nw01769 = ~(nw01768 | nw00564);
  assign nw01770 = nw00575 ? nw01756 : nw01769;
  assign nw01771 = ~\nw05423 [13];
  assign nw01772 = ~\nr00020 [13];
  assign nw01773 = ~\nr00019 [13];
  assign nw01774 = ~\nr00021 [13];
  assign nw01775 = ~\nw05422 [13];
  assign nw01776 = ~\nr00018 [13];
  assign nw01777 = ~\nr00024 [13];
  assign nw01778 = \nr00015  ? nw01777 : nw01776;
  assign nw01779 = nw01375 ? nw01775 : nw01778;
  assign nw01780 = nw01377 ? nw01774 : nw01779;
  assign nw01781 = nw01379 ? nw01773 : nw01780;
  assign nw01782 = nw01381 ? nw01772 : nw01781;
  assign nw01783 = nw01383 ? nw01771 : nw01782;
  assign nw01784 = nw01783 | nw01385;
  assign nw01785 = ~(nw01784 | nw01387);
  assign nw00069 = nw00587 ? nw01770 : nw01785;
  assign nw01786 = ~\nr00064 [14];
  assign nw01787 = ~\nr00064 [30];
  assign nw01788 = address_ext_o[1] ? nw01787 : nw01786;
  assign nw01789 = ~nw01788;
  assign nw01790 = ~\nr00026 [14];
  assign nw01791 = ~\nr00066 [14];
  assign nw01792 = nw00465 ? nw01790 : nw01791;
  assign nw01793 = nw00475 ? nw01591 : nw01792;
  assign nw01794 = nw00484 ? nw01590 : nw01793;
  assign nw01795 = nw00493 ? nw00978 : nw01794;
  assign nw01796 = nw00502 ? nw01589 : nw01795;
  assign nw01797 = nw00510 ? nw01788 : nw01796;
  assign nw01798 = nw00519 ? nw01786 : nw01797;
  assign nw01799 = nw01798 | nw00531;
  assign nw01800 = nw01799 | nw00542;
  assign nw01801 = nw01800 | nw00553;
  assign nw01802 = ~(nw01801 | nw00564);
  assign nw01803 = nw00575 ? nw01789 : nw01802;
  assign nw01804 = ~\nw05423 [14];
  assign nw01805 = ~\nr00020 [14];
  assign nw01806 = ~\nr00019 [14];
  assign nw01807 = ~\nr00021 [14];
  assign nw01808 = ~\nw05422 [14];
  assign nw01809 = ~\nr00018 [14];
  assign nw01810 = ~\nr00024 [14];
  assign nw01811 = \nr00015  ? nw01810 : nw01809;
  assign nw01812 = nw01375 ? nw01808 : nw01811;
  assign nw01813 = nw01377 ? nw01807 : nw01812;
  assign nw01814 = nw01379 ? nw01806 : nw01813;
  assign nw01815 = nw01381 ? nw01805 : nw01814;
  assign nw01816 = nw01383 ? nw01804 : nw01815;
  assign nw01817 = nw01816 | nw01385;
  assign nw01818 = ~(nw01817 | nw01387);
  assign nw00070 = nw00587 ? nw01803 : nw01818;
  assign nw01819 = address_ext_o[1] ? nw00978 : nw01591;
  assign nw01820 = ~nw01819;
  assign nw01821 = ~\nr00026 [15];
  assign nw01822 = ~\nr00066 [15];
  assign nw01823 = nw00465 ? nw01821 : nw01822;
  assign nw01824 = nw00475 ? nw01591 : nw01823;
  assign nw01825 = nw00484 ? nw01590 : nw01824;
  assign nw01826 = nw00493 ? nw00978 : nw01825;
  assign nw01827 = nw00502 ? nw01589 : nw01826;
  assign nw01828 = nw00510 ? nw01819 : nw01827;
  assign nw01829 = nw00519 ? nw01591 : nw01828;
  assign nw01830 = nw01829 | nw00531;
  assign nw01831 = nw01830 | nw00542;
  assign nw01832 = nw01831 | nw00553;
  assign nw01833 = ~(nw01832 | nw00564);
  assign nw01834 = nw00575 ? nw01820 : nw01833;
  assign nw01835 = ~\nw05423 [15];
  assign nw01836 = ~\nr00020 [15];
  assign nw01837 = ~\nr00019 [15];
  assign nw01838 = ~\nr00021 [15];
  assign nw01839 = ~\nw05422 [15];
  assign nw01840 = ~\nr00018 [15];
  assign nw01841 = ~\nr00024 [15];
  assign nw01842 = \nr00015  ? nw01841 : nw01840;
  assign nw01843 = nw01375 ? nw01839 : nw01842;
  assign nw01844 = nw01377 ? nw01838 : nw01843;
  assign nw01845 = nw01379 ? nw01837 : nw01844;
  assign nw01846 = nw01381 ? nw01836 : nw01845;
  assign nw01847 = nw01383 ? nw01835 : nw01846;
  assign nw01848 = nw01847 | nw01385;
  assign nw01849 = ~(nw01848 | nw01387);
  assign nw00071 = nw00587 ? nw01834 : nw01849;
  assign nw01850 = ~\nr00064 [16];
  assign nw01851 = ~\nr00026 [16];
  assign nw01852 = ~\nr00066 [16];
  assign nw01853 = nw00465 ? nw01851 : nw01852;
  assign nw01854 = nw00475 ? nw01591 : nw01853;
  assign nw01855 = nw00484 ? nw01590 : nw01854;
  assign nw01856 = nw00493 ? nw00978 : nw01855;
  assign nw01857 = nw00502 ? nw01589 : nw01856;
  assign nw01858 = nw00510 ? nw01819 : nw01857;
  assign nw01859 = nw00519 ? nw01850 : nw01858;
  assign nw01860 = nw01859 | nw00531;
  assign nw01861 = nw01860 | nw00542;
  assign nw01862 = nw01861 | nw00553;
  assign nw01863 = nw01862 | nw00564;
  assign nw01864 = ~(nw01863 | nw00575);
  assign nw01865 = ~\nw05423 [16];
  assign nw01866 = ~\nr00020 [16];
  assign nw01867 = ~\nr00019 [16];
  assign nw01868 = ~\nr00021 [16];
  assign nw01869 = ~\nw05422 [16];
  assign nw01870 = ~\nr00018 [16];
  assign nw01871 = ~\nr00024 [16];
  assign nw01872 = \nr00015  ? nw01871 : nw01870;
  assign nw01873 = nw01375 ? nw01869 : nw01872;
  assign nw01874 = nw01377 ? nw01868 : nw01873;
  assign nw01875 = nw01379 ? nw01867 : nw01874;
  assign nw01876 = nw01381 ? nw01866 : nw01875;
  assign nw01877 = nw01383 ? nw01865 : nw01876;
  assign nw01878 = nw01877 | nw01385;
  assign nw01879 = ~(nw01878 | nw01387);
  assign nw00072 = nw00587 ? nw01864 : nw01879;
  assign nw01880 = ~\nr00064 [17];
  assign nw01881 = ~\nr00026 [17];
  assign nw01882 = ~\nr00066 [17];
  assign nw01883 = nw00465 ? nw01881 : nw01882;
  assign nw01884 = nw00475 ? nw01591 : nw01883;
  assign nw01885 = nw00484 ? nw01590 : nw01884;
  assign nw01886 = nw00493 ? nw00978 : nw01885;
  assign nw01887 = nw00502 ? nw01589 : nw01886;
  assign nw01888 = nw00510 ? nw01819 : nw01887;
  assign nw01889 = nw00519 ? nw01880 : nw01888;
  assign nw01890 = nw01889 | nw00531;
  assign nw01891 = nw01890 | nw00542;
  assign nw01892 = nw01891 | nw00553;
  assign nw01893 = nw01892 | nw00564;
  assign nw01894 = ~(nw01893 | nw00575);
  assign nw01895 = ~\nw05423 [17];
  assign nw01896 = ~\nr00020 [17];
  assign nw01897 = ~\nr00019 [17];
  assign nw01898 = ~\nr00021 [17];
  assign nw01899 = ~\nw05422 [17];
  assign nw01900 = ~\nr00018 [17];
  assign nw01901 = ~\nr00024 [17];
  assign nw01902 = \nr00015  ? nw01901 : nw01900;
  assign nw01903 = nw01375 ? nw01899 : nw01902;
  assign nw01904 = nw01377 ? nw01898 : nw01903;
  assign nw01905 = nw01379 ? nw01897 : nw01904;
  assign nw01906 = nw01381 ? nw01896 : nw01905;
  assign nw01907 = nw01383 ? nw01895 : nw01906;
  assign nw01908 = nw01907 | nw01385;
  assign nw01909 = ~(nw01908 | nw01387);
  assign nw00073 = nw00587 ? nw01894 : nw01909;
  assign nw01910 = ~\nr00064 [18];
  assign nw01911 = ~\nr00026 [18];
  assign nw01912 = ~\nr00066 [18];
  assign nw01913 = nw00465 ? nw01911 : nw01912;
  assign nw01914 = nw00475 ? nw01591 : nw01913;
  assign nw01915 = nw00484 ? nw01590 : nw01914;
  assign nw01916 = nw00493 ? nw00978 : nw01915;
  assign nw01917 = nw00502 ? nw01589 : nw01916;
  assign nw01918 = nw00510 ? nw01819 : nw01917;
  assign nw01919 = nw00519 ? nw01910 : nw01918;
  assign nw01920 = nw01919 | nw00531;
  assign nw01921 = nw01920 | nw00542;
  assign nw01922 = nw01921 | nw00553;
  assign nw01923 = nw01922 | nw00564;
  assign nw01924 = ~(nw01923 | nw00575);
  assign nw01925 = ~\nw05423 [18];
  assign nw01926 = ~\nr00020 [18];
  assign nw01927 = ~\nr00019 [18];
  assign nw01928 = ~\nr00021 [18];
  assign nw01929 = ~\nw05422 [18];
  assign nw01930 = ~\nr00018 [18];
  assign nw01931 = ~\nr00024 [18];
  assign nw01932 = \nr00015  ? nw01931 : nw01930;
  assign nw01933 = nw01375 ? nw01929 : nw01932;
  assign nw01934 = nw01377 ? nw01928 : nw01933;
  assign nw01935 = nw01379 ? nw01927 : nw01934;
  assign nw01936 = nw01381 ? nw01926 : nw01935;
  assign nw01937 = nw01383 ? nw01925 : nw01936;
  assign nw01938 = nw01937 | nw01385;
  assign nw01939 = ~(nw01938 | nw01387);
  assign nw00074 = nw00587 ? nw01924 : nw01939;
  assign nw01940 = ~\nr00064 [19];
  assign nw01941 = ~\nr00026 [19];
  assign nw01942 = ~\nr00066 [19];
  assign nw01943 = nw00465 ? nw01941 : nw01942;
  assign nw01944 = nw00475 ? nw01591 : nw01943;
  assign nw01945 = nw00484 ? nw01590 : nw01944;
  assign nw01946 = nw00493 ? nw00978 : nw01945;
  assign nw01947 = nw00502 ? nw01589 : nw01946;
  assign nw01948 = nw00510 ? nw01819 : nw01947;
  assign nw01949 = nw00519 ? nw01940 : nw01948;
  assign nw01950 = nw01949 | nw00531;
  assign nw01951 = nw01950 | nw00542;
  assign nw01952 = nw01951 | nw00553;
  assign nw01953 = nw01952 | nw00564;
  assign nw01954 = ~(nw01953 | nw00575);
  assign nw01955 = ~\nw05423 [19];
  assign nw01956 = ~\nr00020 [19];
  assign nw01957 = ~\nr00019 [19];
  assign nw01958 = ~\nr00021 [19];
  assign nw01959 = ~\nw05422 [19];
  assign nw01960 = ~\nr00018 [19];
  assign nw01961 = ~\nr00024 [19];
  assign nw01962 = \nr00015  ? nw01961 : nw01960;
  assign nw01963 = nw01375 ? nw01959 : nw01962;
  assign nw01964 = nw01377 ? nw01958 : nw01963;
  assign nw01965 = nw01379 ? nw01957 : nw01964;
  assign nw01966 = nw01381 ? nw01956 : nw01965;
  assign nw01967 = nw01383 ? nw01955 : nw01966;
  assign nw01968 = nw01967 | nw01385;
  assign nw01969 = ~(nw01968 | nw01387);
  assign nw00075 = nw00587 ? nw01954 : nw01969;
  assign nw01970 = ~\nr00064 [20];
  assign nw01971 = ~\nr00026 [20];
  assign nw01972 = ~\nr00066 [20];
  assign nw01973 = nw00465 ? nw01971 : nw01972;
  assign nw01974 = nw00475 ? nw01591 : nw01973;
  assign nw01975 = nw00484 ? nw01590 : nw01974;
  assign nw01976 = nw00493 ? nw00978 : nw01975;
  assign nw01977 = nw00502 ? nw01589 : nw01976;
  assign nw01978 = nw00510 ? nw01819 : nw01977;
  assign nw01979 = nw00519 ? nw01970 : nw01978;
  assign nw01980 = nw01979 | nw00531;
  assign nw01981 = nw01980 | nw00542;
  assign nw01982 = nw01981 | nw00553;
  assign nw01983 = nw01982 | nw00564;
  assign nw01984 = ~(nw01983 | nw00575);
  assign nw01985 = ~\nw05423 [20];
  assign nw01986 = ~\nr00020 [20];
  assign nw01987 = ~\nr00019 [20];
  assign nw01988 = ~\nr00021 [20];
  assign nw01989 = ~\nw05422 [20];
  assign nw01990 = ~\nr00018 [20];
  assign nw01991 = ~\nr00024 [20];
  assign nw01992 = \nr00015  ? nw01991 : nw01990;
  assign nw01993 = nw01375 ? nw01989 : nw01992;
  assign nw01994 = nw01377 ? nw01988 : nw01993;
  assign nw01995 = nw01379 ? nw01987 : nw01994;
  assign nw01996 = nw01381 ? nw01986 : nw01995;
  assign nw01997 = nw01383 ? nw01985 : nw01996;
  assign nw01998 = nw01997 | nw01385;
  assign nw01999 = ~(nw01998 | nw01387);
  assign nw00077 = nw00587 ? nw01984 : nw01999;
  assign nw02000 = ~\nr00064 [21];
  assign nw02001 = ~\nr00026 [21];
  assign nw02002 = ~\nr00066 [21];
  assign nw02003 = nw00465 ? nw02001 : nw02002;
  assign nw02004 = nw00475 ? nw01591 : nw02003;
  assign nw02005 = nw00484 ? nw01590 : nw02004;
  assign nw02006 = nw00493 ? nw00978 : nw02005;
  assign nw02007 = nw00502 ? nw01589 : nw02006;
  assign nw02008 = nw00510 ? nw01819 : nw02007;
  assign nw02009 = nw00519 ? nw02000 : nw02008;
  assign nw02010 = nw02009 | nw00531;
  assign nw02011 = nw02010 | nw00542;
  assign nw02012 = nw02011 | nw00553;
  assign nw02013 = nw02012 | nw00564;
  assign nw02014 = ~(nw02013 | nw00575);
  assign nw02015 = ~\nw05423 [21];
  assign nw02016 = ~\nr00020 [21];
  assign nw02017 = ~\nr00019 [21];
  assign nw02018 = ~\nr00021 [21];
  assign nw02019 = ~\nw05422 [21];
  assign nw02020 = ~\nr00018 [21];
  assign nw02021 = ~\nr00024 [21];
  assign nw02022 = \nr00015  ? nw02021 : nw02020;
  assign nw02023 = nw01375 ? nw02019 : nw02022;
  assign nw02024 = nw01377 ? nw02018 : nw02023;
  assign nw02025 = nw01379 ? nw02017 : nw02024;
  assign nw02026 = nw01381 ? nw02016 : nw02025;
  assign nw02027 = nw01383 ? nw02015 : nw02026;
  assign nw02028 = nw02027 | nw01385;
  assign nw02029 = ~(nw02028 | nw01387);
  assign nw00078 = nw00587 ? nw02014 : nw02029;
  assign nw02030 = ~\nr00064 [22];
  assign nw02031 = ~\nr00026 [22];
  assign nw02032 = ~\nr00066 [22];
  assign nw02033 = nw00465 ? nw02031 : nw02032;
  assign nw02034 = nw00475 ? nw01591 : nw02033;
  assign nw02035 = nw00484 ? nw01590 : nw02034;
  assign nw02036 = nw00493 ? nw00978 : nw02035;
  assign nw02037 = nw00502 ? nw01589 : nw02036;
  assign nw02038 = nw00510 ? nw01819 : nw02037;
  assign nw02039 = nw00519 ? nw02030 : nw02038;
  assign nw02040 = nw02039 | nw00531;
  assign nw02041 = nw02040 | nw00542;
  assign nw02042 = nw02041 | nw00553;
  assign nw02043 = nw02042 | nw00564;
  assign nw02044 = ~(nw02043 | nw00575);
  assign nw02045 = ~\nw05423 [22];
  assign nw02046 = ~\nr00020 [22];
  assign nw02047 = ~\nr00019 [22];
  assign nw02048 = ~\nr00021 [22];
  assign nw02049 = ~\nw05422 [22];
  assign nw02050 = ~\nr00018 [22];
  assign nw02051 = ~\nr00024 [22];
  assign nw02052 = \nr00015  ? nw02051 : nw02050;
  assign nw02053 = nw01375 ? nw02049 : nw02052;
  assign nw02054 = nw01377 ? nw02048 : nw02053;
  assign nw02055 = nw01379 ? nw02047 : nw02054;
  assign nw02056 = nw01381 ? nw02046 : nw02055;
  assign nw02057 = nw01383 ? nw02045 : nw02056;
  assign nw02058 = nw02057 | nw01385;
  assign nw02059 = ~(nw02058 | nw01387);
  assign nw00079 = nw00587 ? nw02044 : nw02059;
  assign nw02060 = ~\nr00026 [23];
  assign nw02061 = ~\nr00066 [23];
  assign nw02062 = nw00465 ? nw02060 : nw02061;
  assign nw02063 = nw00475 ? nw01591 : nw02062;
  assign nw02064 = nw00484 ? nw01590 : nw02063;
  assign nw02065 = nw00493 ? nw00978 : nw02064;
  assign nw02066 = nw00502 ? nw01589 : nw02065;
  assign nw02067 = nw00510 ? nw01819 : nw02066;
  assign nw02068 = nw00519 ? nw01590 : nw02067;
  assign nw02069 = nw02068 | nw00531;
  assign nw02070 = nw02069 | nw00542;
  assign nw02071 = nw02070 | nw00553;
  assign nw02072 = nw02071 | nw00564;
  assign nw02073 = ~(nw02072 | nw00575);
  assign nw02074 = ~\nw05423 [23];
  assign nw02075 = ~\nr00020 [23];
  assign nw02076 = ~\nr00019 [23];
  assign nw02077 = ~\nr00021 [23];
  assign nw02078 = ~\nw05422 [23];
  assign nw02079 = ~\nr00018 [23];
  assign nw02080 = ~\nr00024 [23];
  assign nw02081 = \nr00015  ? nw02080 : nw02079;
  assign nw02082 = nw01375 ? nw02078 : nw02081;
  assign nw02083 = nw01377 ? nw02077 : nw02082;
  assign nw02084 = nw01379 ? nw02076 : nw02083;
  assign nw02085 = nw01381 ? nw02075 : nw02084;
  assign nw02086 = nw01383 ? nw02074 : nw02085;
  assign nw02087 = nw02086 | nw01385;
  assign nw02088 = ~(nw02087 | nw01387);
  assign nw00080 = nw00587 ? nw02073 : nw02088;
  assign nw02089 = ~\nr00026 [24];
  assign nw02090 = ~\nr00066 [24];
  assign nw02091 = nw00465 ? nw02089 : nw02090;
  assign nw02092 = nw00475 ? nw01591 : nw02091;
  assign nw02093 = nw00484 ? nw01590 : nw02092;
  assign nw02094 = nw00493 ? nw00978 : nw02093;
  assign nw02095 = nw00502 ? nw01589 : nw02094;
  assign nw02096 = nw00510 ? nw01819 : nw02095;
  assign nw02097 = nw00519 ? nw01586 : nw02096;
  assign nw02098 = nw02097 | nw00531;
  assign nw02099 = nw02098 | nw00542;
  assign nw02100 = nw02099 | nw00553;
  assign nw02101 = nw02100 | nw00564;
  assign nw02102 = ~(nw02101 | nw00575);
  assign nw02103 = ~\nw05423 [24];
  assign nw02104 = ~\nr00020 [24];
  assign nw02105 = ~\nr00019 [24];
  assign nw02106 = ~\nr00021 [24];
  assign nw02107 = ~\nw05422 [24];
  assign nw02108 = ~\nr00018 [24];
  assign nw02109 = ~\nr00024 [24];
  assign nw02110 = \nr00015  ? nw02109 : nw02108;
  assign nw02111 = nw01375 ? nw02107 : nw02110;
  assign nw02112 = nw01377 ? nw02106 : nw02111;
  assign nw02113 = nw01379 ? nw02105 : nw02112;
  assign nw02114 = nw01381 ? nw02104 : nw02113;
  assign nw02115 = nw01383 ? nw02103 : nw02114;
  assign nw02116 = nw02115 | nw01385;
  assign nw02117 = ~(nw02116 | nw01387);
  assign nw00081 = nw00587 ? nw02102 : nw02117;
  assign nw02118 = ~\nr00026 [25];
  assign nw02119 = ~\nr00066 [25];
  assign nw02120 = nw00465 ? nw02118 : nw02119;
  assign nw02121 = nw00475 ? nw01591 : nw02120;
  assign nw02122 = nw00484 ? nw01590 : nw02121;
  assign nw02123 = nw00493 ? nw00978 : nw02122;
  assign nw02124 = nw00502 ? nw01589 : nw02123;
  assign nw02125 = nw00510 ? nw01819 : nw02124;
  assign nw02126 = nw00519 ? nw01621 : nw02125;
  assign nw02127 = nw02126 | nw00531;
  assign nw02128 = nw02127 | nw00542;
  assign nw02129 = nw02128 | nw00553;
  assign nw02130 = nw02129 | nw00564;
  assign nw02131 = ~(nw02130 | nw00575);
  assign nw02132 = ~\nw05423 [25];
  assign nw02133 = ~\nr00020 [25];
  assign nw02134 = ~\nr00019 [25];
  assign nw02135 = ~\nr00021 [25];
  assign nw02136 = ~\nw05422 [25];
  assign nw02137 = ~\nr00018 [25];
  assign nw02138 = ~\nr00024 [25];
  assign nw02139 = \nr00015  ? nw02138 : nw02137;
  assign nw02140 = nw01375 ? nw02136 : nw02139;
  assign nw02141 = nw01377 ? nw02135 : nw02140;
  assign nw02142 = nw01379 ? nw02134 : nw02141;
  assign nw02143 = nw01381 ? nw02133 : nw02142;
  assign nw02144 = nw01383 ? nw02132 : nw02143;
  assign nw02145 = nw02144 | nw01385;
  assign nw02146 = ~(nw02145 | nw01387);
  assign nw00082 = nw00587 ? nw02131 : nw02146;
  assign nw02147 = ~\nr00026 [26];
  assign nw02148 = ~\nr00066 [26];
  assign nw02149 = nw00465 ? nw02147 : nw02148;
  assign nw02150 = nw00475 ? nw01591 : nw02149;
  assign nw02151 = nw00484 ? nw01590 : nw02150;
  assign nw02152 = nw00493 ? nw00978 : nw02151;
  assign nw02153 = nw00502 ? nw01589 : nw02152;
  assign nw02154 = nw00510 ? nw01819 : nw02153;
  assign nw02155 = nw00519 ? nw01654 : nw02154;
  assign nw02156 = nw02155 | nw00531;
  assign nw02157 = nw02156 | nw00542;
  assign nw02158 = nw02157 | nw00553;
  assign nw02159 = nw02158 | nw00564;
  assign nw02160 = ~(nw02159 | nw00575);
  assign nw02161 = ~\nw05423 [26];
  assign nw02162 = ~\nr00020 [26];
  assign nw02163 = ~\nr00019 [26];
  assign nw02164 = ~\nr00021 [26];
  assign nw02165 = ~\nw05422 [26];
  assign nw02166 = ~\nr00018 [26];
  assign nw02167 = ~\nr00024 [26];
  assign nw02168 = \nr00015  ? nw02167 : nw02166;
  assign nw02169 = nw01375 ? nw02165 : nw02168;
  assign nw02170 = nw01377 ? nw02164 : nw02169;
  assign nw02171 = nw01379 ? nw02163 : nw02170;
  assign nw02172 = nw01381 ? nw02162 : nw02171;
  assign nw02173 = nw01383 ? nw02161 : nw02172;
  assign nw02174 = nw02173 | nw01385;
  assign nw02175 = ~(nw02174 | nw01387);
  assign nw00083 = nw00587 ? nw02160 : nw02175;
  assign nw02176 = ~\nr00026 [27];
  assign nw02177 = ~\nr00066 [27];
  assign nw02178 = nw00465 ? nw02176 : nw02177;
  assign nw02179 = nw00475 ? nw01591 : nw02178;
  assign nw02180 = nw00484 ? nw01590 : nw02179;
  assign nw02181 = nw00493 ? nw00978 : nw02180;
  assign nw02182 = nw00502 ? nw01589 : nw02181;
  assign nw02183 = nw00510 ? nw01819 : nw02182;
  assign nw02184 = nw00519 ? nw01687 : nw02183;
  assign nw02185 = nw02184 | nw00531;
  assign nw02186 = nw02185 | nw00542;
  assign nw02187 = nw02186 | nw00553;
  assign nw02188 = nw02187 | nw00564;
  assign nw02189 = ~(nw02188 | nw00575);
  assign nw02190 = ~\nw05423 [27];
  assign nw02191 = ~\nr00020 [27];
  assign nw02192 = ~\nr00019 [27];
  assign nw02193 = ~\nr00021 [27];
  assign nw02194 = ~\nw05422 [27];
  assign nw02195 = ~\nr00018 [27];
  assign nw02196 = ~\nr00024 [27];
  assign nw02197 = \nr00015  ? nw02196 : nw02195;
  assign nw02198 = nw01375 ? nw02194 : nw02197;
  assign nw02199 = nw01377 ? nw02193 : nw02198;
  assign nw02200 = nw01379 ? nw02192 : nw02199;
  assign nw02201 = nw01381 ? nw02191 : nw02200;
  assign nw02202 = nw01383 ? nw02190 : nw02201;
  assign nw02203 = nw02202 | nw01385;
  assign nw02204 = ~(nw02203 | nw01387);
  assign nw00084 = nw00587 ? nw02189 : nw02204;
  assign nw02205 = ~\nr00026 [28];
  assign nw02206 = ~\nr00066 [28];
  assign nw02207 = nw00465 ? nw02205 : nw02206;
  assign nw02208 = nw00475 ? nw01591 : nw02207;
  assign nw02209 = nw00484 ? nw01590 : nw02208;
  assign nw02210 = nw00493 ? nw00978 : nw02209;
  assign nw02211 = nw00502 ? nw01589 : nw02210;
  assign nw02212 = nw00510 ? nw01819 : nw02211;
  assign nw02213 = nw00519 ? nw01721 : nw02212;
  assign nw02214 = nw02213 | nw00531;
  assign nw02215 = nw02214 | nw00542;
  assign nw02216 = nw02215 | nw00553;
  assign nw02217 = nw02216 | nw00564;
  assign nw02218 = ~(nw02217 | nw00575);
  assign nw02219 = ~\nw05423 [28];
  assign nw02220 = ~\nr00020 [28];
  assign nw02221 = ~\nr00019 [28];
  assign nw02222 = ~\nr00021 [28];
  assign nw02223 = ~\nw05422 [28];
  assign nw02224 = ~\nr00018 [28];
  assign nw02225 = ~\nr00024 [28];
  assign nw02226 = \nr00015  ? nw02225 : nw02224;
  assign nw02227 = nw01375 ? nw02223 : nw02226;
  assign nw02228 = nw01377 ? nw02222 : nw02227;
  assign nw02229 = nw01379 ? nw02221 : nw02228;
  assign nw02230 = nw01381 ? nw02220 : nw02229;
  assign nw02231 = nw01383 ? nw02219 : nw02230;
  assign nw02232 = nw02231 | nw01385;
  assign nw02233 = ~(nw02232 | nw01387);
  assign nw00085 = nw00587 ? nw02218 : nw02233;
  assign nw02234 = ~\nr00026 [29];
  assign nw02235 = ~\nr00066 [29];
  assign nw02236 = nw00465 ? nw02234 : nw02235;
  assign nw02237 = nw00475 ? nw01591 : nw02236;
  assign nw02238 = nw00484 ? nw01590 : nw02237;
  assign nw02239 = nw00493 ? nw00978 : nw02238;
  assign nw02240 = nw00502 ? nw01589 : nw02239;
  assign nw02241 = nw00510 ? nw01819 : nw02240;
  assign nw02242 = nw00519 ? nw01754 : nw02241;
  assign nw02243 = nw02242 | nw00531;
  assign nw02244 = nw02243 | nw00542;
  assign nw02245 = nw02244 | nw00553;
  assign nw02246 = nw02245 | nw00564;
  assign nw02247 = ~(nw02246 | nw00575);
  assign nw02248 = ~\nw05423 [29];
  assign nw02249 = ~\nr00020 [29];
  assign nw02250 = ~\nr00019 [29];
  assign nw02251 = ~\nr00021 [29];
  assign nw02252 = ~\nw05422 [29];
  assign nw02253 = ~\nr00018 [29];
  assign nw02254 = ~\nr00024 [29];
  assign nw02255 = \nr00015  ? nw02254 : nw02253;
  assign nw02256 = nw01375 ? nw02252 : nw02255;
  assign nw02257 = nw01377 ? nw02251 : nw02256;
  assign nw02258 = nw01379 ? nw02250 : nw02257;
  assign nw02259 = nw01381 ? nw02249 : nw02258;
  assign nw02260 = nw01383 ? nw02248 : nw02259;
  assign nw02261 = nw02260 | nw01385;
  assign nw02262 = ~(nw02261 | nw01387);
  assign nw00086 = nw00587 ? nw02247 : nw02262;
  assign nw02263 = ~\nr00026 [30];
  assign nw02264 = ~\nr00066 [30];
  assign nw02265 = nw00465 ? nw02263 : nw02264;
  assign nw02266 = nw00475 ? nw01591 : nw02265;
  assign nw02267 = nw00484 ? nw01590 : nw02266;
  assign nw02268 = nw00493 ? nw00978 : nw02267;
  assign nw02269 = nw00502 ? nw01589 : nw02268;
  assign nw02270 = nw00510 ? nw01819 : nw02269;
  assign nw02271 = nw00519 ? nw01787 : nw02270;
  assign nw02272 = nw02271 | nw00531;
  assign nw02273 = nw02272 | nw00542;
  assign nw02274 = nw02273 | nw00553;
  assign nw02275 = nw02274 | nw00564;
  assign nw02276 = ~(nw02275 | nw00575);
  assign nw02277 = ~\nw05423 [30];
  assign nw02278 = ~\nr00020 [30];
  assign nw02279 = ~\nr00019 [30];
  assign nw02280 = ~\nr00021 [30];
  assign nw02281 = ~\nw05422 [30];
  assign nw02282 = ~\nr00018 [30];
  assign nw02283 = ~\nr00024 [30];
  assign nw02284 = \nr00015  ? nw02283 : nw02282;
  assign nw02285 = nw01375 ? nw02281 : nw02284;
  assign nw02286 = nw01377 ? nw02280 : nw02285;
  assign nw02287 = nw01379 ? nw02279 : nw02286;
  assign nw02288 = nw01381 ? nw02278 : nw02287;
  assign nw02289 = nw01383 ? nw02277 : nw02288;
  assign nw02290 = nw02289 | nw01385;
  assign nw02291 = ~(nw02290 | nw01387);
  assign nw00088 = nw00587 ? nw02276 : nw02291;
  assign nw02292 = ~\nr00026 [31];
  assign nw02293 = ~\nr00066 [31];
  assign nw02294 = nw00465 ? nw02292 : nw02293;
  assign nw02295 = nw00475 ? nw01591 : nw02294;
  assign nw02296 = nw00484 ? nw01590 : nw02295;
  assign nw02297 = nw00493 ? nw00978 : nw02296;
  assign nw02298 = nw00502 ? nw01589 : nw02297;
  assign nw02299 = nw00510 ? nw01819 : nw02298;
  assign nw02300 = nw00519 ? nw00978 : nw02299;
  assign nw02301 = nw02300 | nw00531;
  assign nw02302 = nw02301 | nw00542;
  assign nw02303 = nw02302 | nw00553;
  assign nw02304 = nw02303 | nw00564;
  assign nw02305 = ~(nw02304 | nw00575);
  assign nw02306 = ~\nw05423 [31];
  assign nw02307 = ~\nr00020 [31];
  assign nw02308 = ~\nr00019 [31];
  assign nw02309 = ~\nr00021 [31];
  assign nw02310 = ~\nw05422 [31];
  assign nw02311 = ~\nr00018 [31];
  assign nw02312 = ~\nr00024 [31];
  assign nw02313 = \nr00015  ? nw02312 : nw02311;
  assign nw02314 = nw01375 ? nw02310 : nw02313;
  assign nw02315 = nw01377 ? nw02309 : nw02314;
  assign nw02316 = nw01379 ? nw02308 : nw02315;
  assign nw02317 = nw01381 ? nw02307 : nw02316;
  assign nw02318 = nw01383 ? nw02306 : nw02317;
  assign nw02319 = nw02318 | nw01385;
  assign nw02320 = ~(nw02319 | nw01387);
  assign nw00089 = nw00587 ? nw02305 : nw02320;
  assign nw00060 = nw00043 ? \nr00064 [15] : \nr00069 [0];
  assign nw00061 = nw00043 ? \nr00064 [16] : \nr00069 [1];
  assign nw00062 = nw00043 ? \nr00064 [17] : \nr00069 [2];
  assign nw00063 = nw00043 ? \nr00064 [18] : \nr00069 [3];
  assign nw00064 = nw00043 ? \nr00064 [19] : \nr00069 [4];
  assign nw00055 = nw00043 ? \nr00064 [20] : \nr00070 [0];
  assign nw00056 = nw00043 ? \nr00064 [21] : \nr00070 [1];
  assign nw00057 = nw00043 ? \nr00064 [22] : \nr00070 [2];
  assign nw00058 = nw00043 ? \nr00064 [23] : \nr00070 [3];
  assign nw00059 = nw00043 ? \nr00064 [24] : \nr00070 [4];
  assign nw02321 = nr00000[0] ? \nr00071[1] [0] : \nr00071[0] [0];
  assign nw02322 = nr00000[0] ? \nr00071[3] [0] : \nr00071[2] [0];
  assign nw02323 = nr00000[1] ? nw02322 : nw02321;
  assign nw02324 = nr00000[0] ? \nr00071[5] [0] : \nr00071[4] [0];
  assign nw02325 = nr00000[0] ? \nr00071[7] [0] : \nr00071[6] [0];
  assign nw02326 = nr00000[1] ? nw02325 : nw02324;
  assign nw02327 = nr00000[2] ? nw02326 : nw02323;
  assign nw02328 = nr00000[0] ? \nr00071[9] [0] : \nr00071[8] [0];
  assign nw02329 = nr00000[0] ? \nr00071[11] [0] : \nr00071[10] [0];
  assign nw02330 = nr00000[1] ? nw02329 : nw02328;
  assign nw02331 = nr00000[0] ? \nr00071[13] [0] : \nr00071[12] [0];
  assign nw02332 = nr00000[0] ? \nr00071[15] [0] : \nr00071[14] [0];
  assign nw02333 = nr00000[1] ? nw02332 : nw02331;
  assign nw02334 = nr00000[2] ? nw02333 : nw02330;
  assign nw02335 = nr00000[3] ? nw02334 : nw02327;
  assign nw02336 = nr00000[0] ? \nr00071[17] [0] : \nr00071[16] [0];
  assign nw02337 = nr00000[0] ? \nr00071[19] [0] : \nr00071[18] [0];
  assign nw02338 = nr00000[1] ? nw02337 : nw02336;
  assign nw02339 = nr00000[0] ? \nr00071[21] [0] : \nr00071[20] [0];
  assign nw02340 = nr00000[0] ? \nr00071[23] [0] : \nr00071[22] [0];
  assign nw02341 = nr00000[1] ? nw02340 : nw02339;
  assign nw02342 = nr00000[2] ? nw02341 : nw02338;
  assign nw02343 = nr00000[0] ? \nr00071[25] [0] : \nr00071[24] [0];
  assign nw02344 = nr00000[0] ? \nr00071[27] [0] : \nr00071[26] [0];
  assign nw02345 = nr00000[1] ? nw02344 : nw02343;
  assign nw02346 = nr00000[0] ? \nr00071[29] [0] : \nr00071[28] [0];
  assign nw02347 = nr00000[0] ? \nr00071[31] [0] : \nr00071[30] [0];
  assign nw02348 = nr00000[1] ? nw02347 : nw02346;
  assign nw02349 = nr00000[2] ? nw02348 : nw02345;
  assign nw02350 = nr00000[3] ? nw02349 : nw02342;
  assign nw00202 = nr00000[4] ? nw02350 : nw02335;
  assign nw02351 = nr00000[0] ? \nr00071[1] [1] : \nr00071[0] [1];
  assign nw02352 = nr00000[0] ? \nr00071[3] [1] : \nr00071[2] [1];
  assign nw02353 = nr00000[1] ? nw02352 : nw02351;
  assign nw02354 = nr00000[0] ? \nr00071[5] [1] : \nr00071[4] [1];
  assign nw02355 = nr00000[0] ? \nr00071[7] [1] : \nr00071[6] [1];
  assign nw02356 = nr00000[1] ? nw02355 : nw02354;
  assign nw02357 = nr00000[2] ? nw02356 : nw02353;
  assign nw02358 = nr00000[0] ? \nr00071[9] [1] : \nr00071[8] [1];
  assign nw02359 = nr00000[0] ? \nr00071[11] [1] : \nr00071[10] [1];
  assign nw02360 = nr00000[1] ? nw02359 : nw02358;
  assign nw02361 = nr00000[0] ? \nr00071[13] [1] : \nr00071[12] [1];
  assign nw02362 = nr00000[0] ? \nr00071[15] [1] : \nr00071[14] [1];
  assign nw02363 = nr00000[1] ? nw02362 : nw02361;
  assign nw02364 = nr00000[2] ? nw02363 : nw02360;
  assign nw02365 = nr00000[3] ? nw02364 : nw02357;
  assign nw02366 = nr00000[0] ? \nr00071[17] [1] : \nr00071[16] [1];
  assign nw02367 = nr00000[0] ? \nr00071[19] [1] : \nr00071[18] [1];
  assign nw02368 = nr00000[1] ? nw02367 : nw02366;
  assign nw02369 = nr00000[0] ? \nr00071[21] [1] : \nr00071[20] [1];
  assign nw02370 = nr00000[0] ? \nr00071[23] [1] : \nr00071[22] [1];
  assign nw02371 = nr00000[1] ? nw02370 : nw02369;
  assign nw02372 = nr00000[2] ? nw02371 : nw02368;
  assign nw02373 = nr00000[0] ? \nr00071[25] [1] : \nr00071[24] [1];
  assign nw02374 = nr00000[0] ? \nr00071[27] [1] : \nr00071[26] [1];
  assign nw02375 = nr00000[1] ? nw02374 : nw02373;
  assign nw02376 = nr00000[0] ? \nr00071[29] [1] : \nr00071[28] [1];
  assign nw02377 = nr00000[0] ? \nr00071[31] [1] : \nr00071[30] [1];
  assign nw02378 = nr00000[1] ? nw02377 : nw02376;
  assign nw02379 = nr00000[2] ? nw02378 : nw02375;
  assign nw02380 = nr00000[3] ? nw02379 : nw02372;
  assign nw00213 = nr00000[4] ? nw02380 : nw02365;
  assign nw02381 = nr00000[0] ? \nr00071[1] [2] : \nr00071[0] [2];
  assign nw02382 = nr00000[0] ? \nr00071[3] [2] : \nr00071[2] [2];
  assign nw02383 = nr00000[1] ? nw02382 : nw02381;
  assign nw02384 = nr00000[0] ? \nr00071[5] [2] : \nr00071[4] [2];
  assign nw02385 = nr00000[0] ? \nr00071[7] [2] : \nr00071[6] [2];
  assign nw02386 = nr00000[1] ? nw02385 : nw02384;
  assign nw02387 = nr00000[2] ? nw02386 : nw02383;
  assign nw02388 = nr00000[0] ? \nr00071[9] [2] : \nr00071[8] [2];
  assign nw02389 = nr00000[0] ? \nr00071[11] [2] : \nr00071[10] [2];
  assign nw02390 = nr00000[1] ? nw02389 : nw02388;
  assign nw02391 = nr00000[0] ? \nr00071[13] [2] : \nr00071[12] [2];
  assign nw02392 = nr00000[0] ? \nr00071[15] [2] : \nr00071[14] [2];
  assign nw02393 = nr00000[1] ? nw02392 : nw02391;
  assign nw02394 = nr00000[2] ? nw02393 : nw02390;
  assign nw02395 = nr00000[3] ? nw02394 : nw02387;
  assign nw02396 = nr00000[0] ? \nr00071[17] [2] : \nr00071[16] [2];
  assign nw02397 = nr00000[0] ? \nr00071[19] [2] : \nr00071[18] [2];
  assign nw02398 = nr00000[1] ? nw02397 : nw02396;
  assign nw02399 = nr00000[0] ? \nr00071[21] [2] : \nr00071[20] [2];
  assign nw02400 = nr00000[0] ? \nr00071[23] [2] : \nr00071[22] [2];
  assign nw02401 = nr00000[1] ? nw02400 : nw02399;
  assign nw02402 = nr00000[2] ? nw02401 : nw02398;
  assign nw02403 = nr00000[0] ? \nr00071[25] [2] : \nr00071[24] [2];
  assign nw02404 = nr00000[0] ? \nr00071[27] [2] : \nr00071[26] [2];
  assign nw02405 = nr00000[1] ? nw02404 : nw02403;
  assign nw02406 = nr00000[0] ? \nr00071[29] [2] : \nr00071[28] [2];
  assign nw02407 = nr00000[0] ? \nr00071[31] [2] : \nr00071[30] [2];
  assign nw02408 = nr00000[1] ? nw02407 : nw02406;
  assign nw02409 = nr00000[2] ? nw02408 : nw02405;
  assign nw02410 = nr00000[3] ? nw02409 : nw02402;
  assign nw00224 = nr00000[4] ? nw02410 : nw02395;
  assign nw02411 = nr00000[0] ? \nr00071[1] [3] : \nr00071[0] [3];
  assign nw02412 = nr00000[0] ? \nr00071[3] [3] : \nr00071[2] [3];
  assign nw02413 = nr00000[1] ? nw02412 : nw02411;
  assign nw02414 = nr00000[0] ? \nr00071[5] [3] : \nr00071[4] [3];
  assign nw02415 = nr00000[0] ? \nr00071[7] [3] : \nr00071[6] [3];
  assign nw02416 = nr00000[1] ? nw02415 : nw02414;
  assign nw02417 = nr00000[2] ? nw02416 : nw02413;
  assign nw02418 = nr00000[0] ? \nr00071[9] [3] : \nr00071[8] [3];
  assign nw02419 = nr00000[0] ? \nr00071[11] [3] : \nr00071[10] [3];
  assign nw02420 = nr00000[1] ? nw02419 : nw02418;
  assign nw02421 = nr00000[0] ? \nr00071[13] [3] : \nr00071[12] [3];
  assign nw02422 = nr00000[0] ? \nr00071[15] [3] : \nr00071[14] [3];
  assign nw02423 = nr00000[1] ? nw02422 : nw02421;
  assign nw02424 = nr00000[2] ? nw02423 : nw02420;
  assign nw02425 = nr00000[3] ? nw02424 : nw02417;
  assign nw02426 = nr00000[0] ? \nr00071[17] [3] : \nr00071[16] [3];
  assign nw02427 = nr00000[0] ? \nr00071[19] [3] : \nr00071[18] [3];
  assign nw02428 = nr00000[1] ? nw02427 : nw02426;
  assign nw02429 = nr00000[0] ? \nr00071[21] [3] : \nr00071[20] [3];
  assign nw02430 = nr00000[0] ? \nr00071[23] [3] : \nr00071[22] [3];
  assign nw02431 = nr00000[1] ? nw02430 : nw02429;
  assign nw02432 = nr00000[2] ? nw02431 : nw02428;
  assign nw02433 = nr00000[0] ? \nr00071[25] [3] : \nr00071[24] [3];
  assign nw02434 = nr00000[0] ? \nr00071[27] [3] : \nr00071[26] [3];
  assign nw02435 = nr00000[1] ? nw02434 : nw02433;
  assign nw02436 = nr00000[0] ? \nr00071[29] [3] : \nr00071[28] [3];
  assign nw02437 = nr00000[0] ? \nr00071[31] [3] : \nr00071[30] [3];
  assign nw02438 = nr00000[1] ? nw02437 : nw02436;
  assign nw02439 = nr00000[2] ? nw02438 : nw02435;
  assign nw02440 = nr00000[3] ? nw02439 : nw02432;
  assign nw00227 = nr00000[4] ? nw02440 : nw02425;
  assign nw02441 = nr00000[0] ? \nr00071[1] [4] : \nr00071[0] [4];
  assign nw02442 = nr00000[0] ? \nr00071[3] [4] : \nr00071[2] [4];
  assign nw02443 = nr00000[1] ? nw02442 : nw02441;
  assign nw02444 = nr00000[0] ? \nr00071[5] [4] : \nr00071[4] [4];
  assign nw02445 = nr00000[0] ? \nr00071[7] [4] : \nr00071[6] [4];
  assign nw02446 = nr00000[1] ? nw02445 : nw02444;
  assign nw02447 = nr00000[2] ? nw02446 : nw02443;
  assign nw02448 = nr00000[0] ? \nr00071[9] [4] : \nr00071[8] [4];
  assign nw02449 = nr00000[0] ? \nr00071[11] [4] : \nr00071[10] [4];
  assign nw02450 = nr00000[1] ? nw02449 : nw02448;
  assign nw02451 = nr00000[0] ? \nr00071[13] [4] : \nr00071[12] [4];
  assign nw02452 = nr00000[0] ? \nr00071[15] [4] : \nr00071[14] [4];
  assign nw02453 = nr00000[1] ? nw02452 : nw02451;
  assign nw02454 = nr00000[2] ? nw02453 : nw02450;
  assign nw02455 = nr00000[3] ? nw02454 : nw02447;
  assign nw02456 = nr00000[0] ? \nr00071[17] [4] : \nr00071[16] [4];
  assign nw02457 = nr00000[0] ? \nr00071[19] [4] : \nr00071[18] [4];
  assign nw02458 = nr00000[1] ? nw02457 : nw02456;
  assign nw02459 = nr00000[0] ? \nr00071[21] [4] : \nr00071[20] [4];
  assign nw02460 = nr00000[0] ? \nr00071[23] [4] : \nr00071[22] [4];
  assign nw02461 = nr00000[1] ? nw02460 : nw02459;
  assign nw02462 = nr00000[2] ? nw02461 : nw02458;
  assign nw02463 = nr00000[0] ? \nr00071[25] [4] : \nr00071[24] [4];
  assign nw02464 = nr00000[0] ? \nr00071[27] [4] : \nr00071[26] [4];
  assign nw02465 = nr00000[1] ? nw02464 : nw02463;
  assign nw02466 = nr00000[0] ? \nr00071[29] [4] : \nr00071[28] [4];
  assign nw02467 = nr00000[0] ? \nr00071[31] [4] : \nr00071[30] [4];
  assign nw02468 = nr00000[1] ? nw02467 : nw02466;
  assign nw02469 = nr00000[2] ? nw02468 : nw02465;
  assign nw02470 = nr00000[3] ? nw02469 : nw02462;
  assign nw00228 = nr00000[4] ? nw02470 : nw02455;
  assign nw02471 = nr00000[0] ? \nr00071[1] [5] : \nr00071[0] [5];
  assign nw02472 = nr00000[0] ? \nr00071[3] [5] : \nr00071[2] [5];
  assign nw02473 = nr00000[1] ? nw02472 : nw02471;
  assign nw02474 = nr00000[0] ? \nr00071[5] [5] : \nr00071[4] [5];
  assign nw02475 = nr00000[0] ? \nr00071[7] [5] : \nr00071[6] [5];
  assign nw02476 = nr00000[1] ? nw02475 : nw02474;
  assign nw02477 = nr00000[2] ? nw02476 : nw02473;
  assign nw02478 = nr00000[0] ? \nr00071[9] [5] : \nr00071[8] [5];
  assign nw02479 = nr00000[0] ? \nr00071[11] [5] : \nr00071[10] [5];
  assign nw02480 = nr00000[1] ? nw02479 : nw02478;
  assign nw02481 = nr00000[0] ? \nr00071[13] [5] : \nr00071[12] [5];
  assign nw02482 = nr00000[0] ? \nr00071[15] [5] : \nr00071[14] [5];
  assign nw02483 = nr00000[1] ? nw02482 : nw02481;
  assign nw02484 = nr00000[2] ? nw02483 : nw02480;
  assign nw02485 = nr00000[3] ? nw02484 : nw02477;
  assign nw02486 = nr00000[0] ? \nr00071[17] [5] : \nr00071[16] [5];
  assign nw02487 = nr00000[0] ? \nr00071[19] [5] : \nr00071[18] [5];
  assign nw02488 = nr00000[1] ? nw02487 : nw02486;
  assign nw02489 = nr00000[0] ? \nr00071[21] [5] : \nr00071[20] [5];
  assign nw02490 = nr00000[0] ? \nr00071[23] [5] : \nr00071[22] [5];
  assign nw02491 = nr00000[1] ? nw02490 : nw02489;
  assign nw02492 = nr00000[2] ? nw02491 : nw02488;
  assign nw02493 = nr00000[0] ? \nr00071[25] [5] : \nr00071[24] [5];
  assign nw02494 = nr00000[0] ? \nr00071[27] [5] : \nr00071[26] [5];
  assign nw02495 = nr00000[1] ? nw02494 : nw02493;
  assign nw02496 = nr00000[0] ? \nr00071[29] [5] : \nr00071[28] [5];
  assign nw02497 = nr00000[0] ? \nr00071[31] [5] : \nr00071[30] [5];
  assign nw02498 = nr00000[1] ? nw02497 : nw02496;
  assign nw02499 = nr00000[2] ? nw02498 : nw02495;
  assign nw02500 = nr00000[3] ? nw02499 : nw02492;
  assign nw00229 = nr00000[4] ? nw02500 : nw02485;
  assign nw02501 = nr00000[0] ? \nr00071[1] [6] : \nr00071[0] [6];
  assign nw02502 = nr00000[0] ? \nr00071[3] [6] : \nr00071[2] [6];
  assign nw02503 = nr00000[1] ? nw02502 : nw02501;
  assign nw02504 = nr00000[0] ? \nr00071[5] [6] : \nr00071[4] [6];
  assign nw02505 = nr00000[0] ? \nr00071[7] [6] : \nr00071[6] [6];
  assign nw02506 = nr00000[1] ? nw02505 : nw02504;
  assign nw02507 = nr00000[2] ? nw02506 : nw02503;
  assign nw02508 = nr00000[0] ? \nr00071[9] [6] : \nr00071[8] [6];
  assign nw02509 = nr00000[0] ? \nr00071[11] [6] : \nr00071[10] [6];
  assign nw02510 = nr00000[1] ? nw02509 : nw02508;
  assign nw02511 = nr00000[0] ? \nr00071[13] [6] : \nr00071[12] [6];
  assign nw02512 = nr00000[0] ? \nr00071[15] [6] : \nr00071[14] [6];
  assign nw02513 = nr00000[1] ? nw02512 : nw02511;
  assign nw02514 = nr00000[2] ? nw02513 : nw02510;
  assign nw02515 = nr00000[3] ? nw02514 : nw02507;
  assign nw02516 = nr00000[0] ? \nr00071[17] [6] : \nr00071[16] [6];
  assign nw02517 = nr00000[0] ? \nr00071[19] [6] : \nr00071[18] [6];
  assign nw02518 = nr00000[1] ? nw02517 : nw02516;
  assign nw02519 = nr00000[0] ? \nr00071[21] [6] : \nr00071[20] [6];
  assign nw02520 = nr00000[0] ? \nr00071[23] [6] : \nr00071[22] [6];
  assign nw02521 = nr00000[1] ? nw02520 : nw02519;
  assign nw02522 = nr00000[2] ? nw02521 : nw02518;
  assign nw02523 = nr00000[0] ? \nr00071[25] [6] : \nr00071[24] [6];
  assign nw02524 = nr00000[0] ? \nr00071[27] [6] : \nr00071[26] [6];
  assign nw02525 = nr00000[1] ? nw02524 : nw02523;
  assign nw02526 = nr00000[0] ? \nr00071[29] [6] : \nr00071[28] [6];
  assign nw02527 = nr00000[0] ? \nr00071[31] [6] : \nr00071[30] [6];
  assign nw02528 = nr00000[1] ? nw02527 : nw02526;
  assign nw02529 = nr00000[2] ? nw02528 : nw02525;
  assign nw02530 = nr00000[3] ? nw02529 : nw02522;
  assign nw00230 = nr00000[4] ? nw02530 : nw02515;
  assign nw02531 = nr00000[0] ? \nr00071[1] [7] : \nr00071[0] [7];
  assign nw02532 = nr00000[0] ? \nr00071[3] [7] : \nr00071[2] [7];
  assign nw02533 = nr00000[1] ? nw02532 : nw02531;
  assign nw02534 = nr00000[0] ? \nr00071[5] [7] : \nr00071[4] [7];
  assign nw02535 = nr00000[0] ? \nr00071[7] [7] : \nr00071[6] [7];
  assign nw02536 = nr00000[1] ? nw02535 : nw02534;
  assign nw02537 = nr00000[2] ? nw02536 : nw02533;
  assign nw02538 = nr00000[0] ? \nr00071[9] [7] : \nr00071[8] [7];
  assign nw02539 = nr00000[0] ? \nr00071[11] [7] : \nr00071[10] [7];
  assign nw02540 = nr00000[1] ? nw02539 : nw02538;
  assign nw02541 = nr00000[0] ? \nr00071[13] [7] : \nr00071[12] [7];
  assign nw02542 = nr00000[0] ? \nr00071[15] [7] : \nr00071[14] [7];
  assign nw02543 = nr00000[1] ? nw02542 : nw02541;
  assign nw02544 = nr00000[2] ? nw02543 : nw02540;
  assign nw02545 = nr00000[3] ? nw02544 : nw02537;
  assign nw02546 = nr00000[0] ? \nr00071[17] [7] : \nr00071[16] [7];
  assign nw02547 = nr00000[0] ? \nr00071[19] [7] : \nr00071[18] [7];
  assign nw02548 = nr00000[1] ? nw02547 : nw02546;
  assign nw02549 = nr00000[0] ? \nr00071[21] [7] : \nr00071[20] [7];
  assign nw02550 = nr00000[0] ? \nr00071[23] [7] : \nr00071[22] [7];
  assign nw02551 = nr00000[1] ? nw02550 : nw02549;
  assign nw02552 = nr00000[2] ? nw02551 : nw02548;
  assign nw02553 = nr00000[0] ? \nr00071[25] [7] : \nr00071[24] [7];
  assign nw02554 = nr00000[0] ? \nr00071[27] [7] : \nr00071[26] [7];
  assign nw02555 = nr00000[1] ? nw02554 : nw02553;
  assign nw02556 = nr00000[0] ? \nr00071[29] [7] : \nr00071[28] [7];
  assign nw02557 = nr00000[0] ? \nr00071[31] [7] : \nr00071[30] [7];
  assign nw02558 = nr00000[1] ? nw02557 : nw02556;
  assign nw02559 = nr00000[2] ? nw02558 : nw02555;
  assign nw02560 = nr00000[3] ? nw02559 : nw02552;
  assign nw00231 = nr00000[4] ? nw02560 : nw02545;
  assign nw02561 = nr00000[0] ? \nr00071[1] [8] : \nr00071[0] [8];
  assign nw02562 = nr00000[0] ? \nr00071[3] [8] : \nr00071[2] [8];
  assign nw02563 = nr00000[1] ? nw02562 : nw02561;
  assign nw02564 = nr00000[0] ? \nr00071[5] [8] : \nr00071[4] [8];
  assign nw02565 = nr00000[0] ? \nr00071[7] [8] : \nr00071[6] [8];
  assign nw02566 = nr00000[1] ? nw02565 : nw02564;
  assign nw02567 = nr00000[2] ? nw02566 : nw02563;
  assign nw02568 = nr00000[0] ? \nr00071[9] [8] : \nr00071[8] [8];
  assign nw02569 = nr00000[0] ? \nr00071[11] [8] : \nr00071[10] [8];
  assign nw02570 = nr00000[1] ? nw02569 : nw02568;
  assign nw02571 = nr00000[0] ? \nr00071[13] [8] : \nr00071[12] [8];
  assign nw02572 = nr00000[0] ? \nr00071[15] [8] : \nr00071[14] [8];
  assign nw02573 = nr00000[1] ? nw02572 : nw02571;
  assign nw02574 = nr00000[2] ? nw02573 : nw02570;
  assign nw02575 = nr00000[3] ? nw02574 : nw02567;
  assign nw02576 = nr00000[0] ? \nr00071[17] [8] : \nr00071[16] [8];
  assign nw02577 = nr00000[0] ? \nr00071[19] [8] : \nr00071[18] [8];
  assign nw02578 = nr00000[1] ? nw02577 : nw02576;
  assign nw02579 = nr00000[0] ? \nr00071[21] [8] : \nr00071[20] [8];
  assign nw02580 = nr00000[0] ? \nr00071[23] [8] : \nr00071[22] [8];
  assign nw02581 = nr00000[1] ? nw02580 : nw02579;
  assign nw02582 = nr00000[2] ? nw02581 : nw02578;
  assign nw02583 = nr00000[0] ? \nr00071[25] [8] : \nr00071[24] [8];
  assign nw02584 = nr00000[0] ? \nr00071[27] [8] : \nr00071[26] [8];
  assign nw02585 = nr00000[1] ? nw02584 : nw02583;
  assign nw02586 = nr00000[0] ? \nr00071[29] [8] : \nr00071[28] [8];
  assign nw02587 = nr00000[0] ? \nr00071[31] [8] : \nr00071[30] [8];
  assign nw02588 = nr00000[1] ? nw02587 : nw02586;
  assign nw02589 = nr00000[2] ? nw02588 : nw02585;
  assign nw02590 = nr00000[3] ? nw02589 : nw02582;
  assign nw00232 = nr00000[4] ? nw02590 : nw02575;
  assign nw02591 = nr00000[0] ? \nr00071[1] [9] : \nr00071[0] [9];
  assign nw02592 = nr00000[0] ? \nr00071[3] [9] : \nr00071[2] [9];
  assign nw02593 = nr00000[1] ? nw02592 : nw02591;
  assign nw02594 = nr00000[0] ? \nr00071[5] [9] : \nr00071[4] [9];
  assign nw02595 = nr00000[0] ? \nr00071[7] [9] : \nr00071[6] [9];
  assign nw02596 = nr00000[1] ? nw02595 : nw02594;
  assign nw02597 = nr00000[2] ? nw02596 : nw02593;
  assign nw02598 = nr00000[0] ? \nr00071[9] [9] : \nr00071[8] [9];
  assign nw02599 = nr00000[0] ? \nr00071[11] [9] : \nr00071[10] [9];
  assign nw02600 = nr00000[1] ? nw02599 : nw02598;
  assign nw02601 = nr00000[0] ? \nr00071[13] [9] : \nr00071[12] [9];
  assign nw02602 = nr00000[0] ? \nr00071[15] [9] : \nr00071[14] [9];
  assign nw02603 = nr00000[1] ? nw02602 : nw02601;
  assign nw02604 = nr00000[2] ? nw02603 : nw02600;
  assign nw02605 = nr00000[3] ? nw02604 : nw02597;
  assign nw02606 = nr00000[0] ? \nr00071[17] [9] : \nr00071[16] [9];
  assign nw02607 = nr00000[0] ? \nr00071[19] [9] : \nr00071[18] [9];
  assign nw02608 = nr00000[1] ? nw02607 : nw02606;
  assign nw02609 = nr00000[0] ? \nr00071[21] [9] : \nr00071[20] [9];
  assign nw02610 = nr00000[0] ? \nr00071[23] [9] : \nr00071[22] [9];
  assign nw02611 = nr00000[1] ? nw02610 : nw02609;
  assign nw02612 = nr00000[2] ? nw02611 : nw02608;
  assign nw02613 = nr00000[0] ? \nr00071[25] [9] : \nr00071[24] [9];
  assign nw02614 = nr00000[0] ? \nr00071[27] [9] : \nr00071[26] [9];
  assign nw02615 = nr00000[1] ? nw02614 : nw02613;
  assign nw02616 = nr00000[0] ? \nr00071[29] [9] : \nr00071[28] [9];
  assign nw02617 = nr00000[0] ? \nr00071[31] [9] : \nr00071[30] [9];
  assign nw02618 = nr00000[1] ? nw02617 : nw02616;
  assign nw02619 = nr00000[2] ? nw02618 : nw02615;
  assign nw02620 = nr00000[3] ? nw02619 : nw02612;
  assign nw00233 = nr00000[4] ? nw02620 : nw02605;
  assign nw02621 = nr00000[0] ? \nr00071[1] [10] : \nr00071[0] [10];
  assign nw02622 = nr00000[0] ? \nr00071[3] [10] : \nr00071[2] [10];
  assign nw02623 = nr00000[1] ? nw02622 : nw02621;
  assign nw02624 = nr00000[0] ? \nr00071[5] [10] : \nr00071[4] [10];
  assign nw02625 = nr00000[0] ? \nr00071[7] [10] : \nr00071[6] [10];
  assign nw02626 = nr00000[1] ? nw02625 : nw02624;
  assign nw02627 = nr00000[2] ? nw02626 : nw02623;
  assign nw02628 = nr00000[0] ? \nr00071[9] [10] : \nr00071[8] [10];
  assign nw02629 = nr00000[0] ? \nr00071[11] [10] : \nr00071[10] [10];
  assign nw02630 = nr00000[1] ? nw02629 : nw02628;
  assign nw02631 = nr00000[0] ? \nr00071[13] [10] : \nr00071[12] [10];
  assign nw02632 = nr00000[0] ? \nr00071[15] [10] : \nr00071[14] [10];
  assign nw02633 = nr00000[1] ? nw02632 : nw02631;
  assign nw02634 = nr00000[2] ? nw02633 : nw02630;
  assign nw02635 = nr00000[3] ? nw02634 : nw02627;
  assign nw02636 = nr00000[0] ? \nr00071[17] [10] : \nr00071[16] [10];
  assign nw02637 = nr00000[0] ? \nr00071[19] [10] : \nr00071[18] [10];
  assign nw02638 = nr00000[1] ? nw02637 : nw02636;
  assign nw02639 = nr00000[0] ? \nr00071[21] [10] : \nr00071[20] [10];
  assign nw02640 = nr00000[0] ? \nr00071[23] [10] : \nr00071[22] [10];
  assign nw02641 = nr00000[1] ? nw02640 : nw02639;
  assign nw02642 = nr00000[2] ? nw02641 : nw02638;
  assign nw02643 = nr00000[0] ? \nr00071[25] [10] : \nr00071[24] [10];
  assign nw02644 = nr00000[0] ? \nr00071[27] [10] : \nr00071[26] [10];
  assign nw02645 = nr00000[1] ? nw02644 : nw02643;
  assign nw02646 = nr00000[0] ? \nr00071[29] [10] : \nr00071[28] [10];
  assign nw02647 = nr00000[0] ? \nr00071[31] [10] : \nr00071[30] [10];
  assign nw02648 = nr00000[1] ? nw02647 : nw02646;
  assign nw02649 = nr00000[2] ? nw02648 : nw02645;
  assign nw02650 = nr00000[3] ? nw02649 : nw02642;
  assign nw00203 = nr00000[4] ? nw02650 : nw02635;
  assign nw02651 = nr00000[0] ? \nr00071[1] [11] : \nr00071[0] [11];
  assign nw02652 = nr00000[0] ? \nr00071[3] [11] : \nr00071[2] [11];
  assign nw02653 = nr00000[1] ? nw02652 : nw02651;
  assign nw02654 = nr00000[0] ? \nr00071[5] [11] : \nr00071[4] [11];
  assign nw02655 = nr00000[0] ? \nr00071[7] [11] : \nr00071[6] [11];
  assign nw02656 = nr00000[1] ? nw02655 : nw02654;
  assign nw02657 = nr00000[2] ? nw02656 : nw02653;
  assign nw02658 = nr00000[0] ? \nr00071[9] [11] : \nr00071[8] [11];
  assign nw02659 = nr00000[0] ? \nr00071[11] [11] : \nr00071[10] [11];
  assign nw02660 = nr00000[1] ? nw02659 : nw02658;
  assign nw02661 = nr00000[0] ? \nr00071[13] [11] : \nr00071[12] [11];
  assign nw02662 = nr00000[0] ? \nr00071[15] [11] : \nr00071[14] [11];
  assign nw02663 = nr00000[1] ? nw02662 : nw02661;
  assign nw02664 = nr00000[2] ? nw02663 : nw02660;
  assign nw02665 = nr00000[3] ? nw02664 : nw02657;
  assign nw02666 = nr00000[0] ? \nr00071[17] [11] : \nr00071[16] [11];
  assign nw02667 = nr00000[0] ? \nr00071[19] [11] : \nr00071[18] [11];
  assign nw02668 = nr00000[1] ? nw02667 : nw02666;
  assign nw02669 = nr00000[0] ? \nr00071[21] [11] : \nr00071[20] [11];
  assign nw02670 = nr00000[0] ? \nr00071[23] [11] : \nr00071[22] [11];
  assign nw02671 = nr00000[1] ? nw02670 : nw02669;
  assign nw02672 = nr00000[2] ? nw02671 : nw02668;
  assign nw02673 = nr00000[0] ? \nr00071[25] [11] : \nr00071[24] [11];
  assign nw02674 = nr00000[0] ? \nr00071[27] [11] : \nr00071[26] [11];
  assign nw02675 = nr00000[1] ? nw02674 : nw02673;
  assign nw02676 = nr00000[0] ? \nr00071[29] [11] : \nr00071[28] [11];
  assign nw02677 = nr00000[0] ? \nr00071[31] [11] : \nr00071[30] [11];
  assign nw02678 = nr00000[1] ? nw02677 : nw02676;
  assign nw02679 = nr00000[2] ? nw02678 : nw02675;
  assign nw02680 = nr00000[3] ? nw02679 : nw02672;
  assign nw00204 = nr00000[4] ? nw02680 : nw02665;
  assign nw02681 = nr00000[0] ? \nr00071[1] [12] : \nr00071[0] [12];
  assign nw02682 = nr00000[0] ? \nr00071[3] [12] : \nr00071[2] [12];
  assign nw02683 = nr00000[1] ? nw02682 : nw02681;
  assign nw02684 = nr00000[0] ? \nr00071[5] [12] : \nr00071[4] [12];
  assign nw02685 = nr00000[0] ? \nr00071[7] [12] : \nr00071[6] [12];
  assign nw02686 = nr00000[1] ? nw02685 : nw02684;
  assign nw02687 = nr00000[2] ? nw02686 : nw02683;
  assign nw02688 = nr00000[0] ? \nr00071[9] [12] : \nr00071[8] [12];
  assign nw02689 = nr00000[0] ? \nr00071[11] [12] : \nr00071[10] [12];
  assign nw02690 = nr00000[1] ? nw02689 : nw02688;
  assign nw02691 = nr00000[0] ? \nr00071[13] [12] : \nr00071[12] [12];
  assign nw02692 = nr00000[0] ? \nr00071[15] [12] : \nr00071[14] [12];
  assign nw02693 = nr00000[1] ? nw02692 : nw02691;
  assign nw02694 = nr00000[2] ? nw02693 : nw02690;
  assign nw02695 = nr00000[3] ? nw02694 : nw02687;
  assign nw02696 = nr00000[0] ? \nr00071[17] [12] : \nr00071[16] [12];
  assign nw02697 = nr00000[0] ? \nr00071[19] [12] : \nr00071[18] [12];
  assign nw02698 = nr00000[1] ? nw02697 : nw02696;
  assign nw02699 = nr00000[0] ? \nr00071[21] [12] : \nr00071[20] [12];
  assign nw02700 = nr00000[0] ? \nr00071[23] [12] : \nr00071[22] [12];
  assign nw02701 = nr00000[1] ? nw02700 : nw02699;
  assign nw02702 = nr00000[2] ? nw02701 : nw02698;
  assign nw02703 = nr00000[0] ? \nr00071[25] [12] : \nr00071[24] [12];
  assign nw02704 = nr00000[0] ? \nr00071[27] [12] : \nr00071[26] [12];
  assign nw02705 = nr00000[1] ? nw02704 : nw02703;
  assign nw02706 = nr00000[0] ? \nr00071[29] [12] : \nr00071[28] [12];
  assign nw02707 = nr00000[0] ? \nr00071[31] [12] : \nr00071[30] [12];
  assign nw02708 = nr00000[1] ? nw02707 : nw02706;
  assign nw02709 = nr00000[2] ? nw02708 : nw02705;
  assign nw02710 = nr00000[3] ? nw02709 : nw02702;
  assign nw00205 = nr00000[4] ? nw02710 : nw02695;
  assign nw02711 = nr00000[0] ? \nr00071[1] [13] : \nr00071[0] [13];
  assign nw02712 = nr00000[0] ? \nr00071[3] [13] : \nr00071[2] [13];
  assign nw02713 = nr00000[1] ? nw02712 : nw02711;
  assign nw02714 = nr00000[0] ? \nr00071[5] [13] : \nr00071[4] [13];
  assign nw02715 = nr00000[0] ? \nr00071[7] [13] : \nr00071[6] [13];
  assign nw02716 = nr00000[1] ? nw02715 : nw02714;
  assign nw02717 = nr00000[2] ? nw02716 : nw02713;
  assign nw02718 = nr00000[0] ? \nr00071[9] [13] : \nr00071[8] [13];
  assign nw02719 = nr00000[0] ? \nr00071[11] [13] : \nr00071[10] [13];
  assign nw02720 = nr00000[1] ? nw02719 : nw02718;
  assign nw02721 = nr00000[0] ? \nr00071[13] [13] : \nr00071[12] [13];
  assign nw02722 = nr00000[0] ? \nr00071[15] [13] : \nr00071[14] [13];
  assign nw02723 = nr00000[1] ? nw02722 : nw02721;
  assign nw02724 = nr00000[2] ? nw02723 : nw02720;
  assign nw02725 = nr00000[3] ? nw02724 : nw02717;
  assign nw02726 = nr00000[0] ? \nr00071[17] [13] : \nr00071[16] [13];
  assign nw02727 = nr00000[0] ? \nr00071[19] [13] : \nr00071[18] [13];
  assign nw02728 = nr00000[1] ? nw02727 : nw02726;
  assign nw02729 = nr00000[0] ? \nr00071[21] [13] : \nr00071[20] [13];
  assign nw02730 = nr00000[0] ? \nr00071[23] [13] : \nr00071[22] [13];
  assign nw02731 = nr00000[1] ? nw02730 : nw02729;
  assign nw02732 = nr00000[2] ? nw02731 : nw02728;
  assign nw02733 = nr00000[0] ? \nr00071[25] [13] : \nr00071[24] [13];
  assign nw02734 = nr00000[0] ? \nr00071[27] [13] : \nr00071[26] [13];
  assign nw02735 = nr00000[1] ? nw02734 : nw02733;
  assign nw02736 = nr00000[0] ? \nr00071[29] [13] : \nr00071[28] [13];
  assign nw02737 = nr00000[0] ? \nr00071[31] [13] : \nr00071[30] [13];
  assign nw02738 = nr00000[1] ? nw02737 : nw02736;
  assign nw02739 = nr00000[2] ? nw02738 : nw02735;
  assign nw02740 = nr00000[3] ? nw02739 : nw02732;
  assign nw00206 = nr00000[4] ? nw02740 : nw02725;
  assign nw02741 = nr00000[0] ? \nr00071[1] [14] : \nr00071[0] [14];
  assign nw02742 = nr00000[0] ? \nr00071[3] [14] : \nr00071[2] [14];
  assign nw02743 = nr00000[1] ? nw02742 : nw02741;
  assign nw02744 = nr00000[0] ? \nr00071[5] [14] : \nr00071[4] [14];
  assign nw02745 = nr00000[0] ? \nr00071[7] [14] : \nr00071[6] [14];
  assign nw02746 = nr00000[1] ? nw02745 : nw02744;
  assign nw02747 = nr00000[2] ? nw02746 : nw02743;
  assign nw02748 = nr00000[0] ? \nr00071[9] [14] : \nr00071[8] [14];
  assign nw02749 = nr00000[0] ? \nr00071[11] [14] : \nr00071[10] [14];
  assign nw02750 = nr00000[1] ? nw02749 : nw02748;
  assign nw02751 = nr00000[0] ? \nr00071[13] [14] : \nr00071[12] [14];
  assign nw02752 = nr00000[0] ? \nr00071[15] [14] : \nr00071[14] [14];
  assign nw02753 = nr00000[1] ? nw02752 : nw02751;
  assign nw02754 = nr00000[2] ? nw02753 : nw02750;
  assign nw02755 = nr00000[3] ? nw02754 : nw02747;
  assign nw02756 = nr00000[0] ? \nr00071[17] [14] : \nr00071[16] [14];
  assign nw02757 = nr00000[0] ? \nr00071[19] [14] : \nr00071[18] [14];
  assign nw02758 = nr00000[1] ? nw02757 : nw02756;
  assign nw02759 = nr00000[0] ? \nr00071[21] [14] : \nr00071[20] [14];
  assign nw02760 = nr00000[0] ? \nr00071[23] [14] : \nr00071[22] [14];
  assign nw02761 = nr00000[1] ? nw02760 : nw02759;
  assign nw02762 = nr00000[2] ? nw02761 : nw02758;
  assign nw02763 = nr00000[0] ? \nr00071[25] [14] : \nr00071[24] [14];
  assign nw02764 = nr00000[0] ? \nr00071[27] [14] : \nr00071[26] [14];
  assign nw02765 = nr00000[1] ? nw02764 : nw02763;
  assign nw02766 = nr00000[0] ? \nr00071[29] [14] : \nr00071[28] [14];
  assign nw02767 = nr00000[0] ? \nr00071[31] [14] : \nr00071[30] [14];
  assign nw02768 = nr00000[1] ? nw02767 : nw02766;
  assign nw02769 = nr00000[2] ? nw02768 : nw02765;
  assign nw02770 = nr00000[3] ? nw02769 : nw02762;
  assign nw00207 = nr00000[4] ? nw02770 : nw02755;
  assign nw02771 = nr00000[0] ? \nr00071[1] [15] : \nr00071[0] [15];
  assign nw02772 = nr00000[0] ? \nr00071[3] [15] : \nr00071[2] [15];
  assign nw02773 = nr00000[1] ? nw02772 : nw02771;
  assign nw02774 = nr00000[0] ? \nr00071[5] [15] : \nr00071[4] [15];
  assign nw02775 = nr00000[0] ? \nr00071[7] [15] : \nr00071[6] [15];
  assign nw02776 = nr00000[1] ? nw02775 : nw02774;
  assign nw02777 = nr00000[2] ? nw02776 : nw02773;
  assign nw02778 = nr00000[0] ? \nr00071[9] [15] : \nr00071[8] [15];
  assign nw02779 = nr00000[0] ? \nr00071[11] [15] : \nr00071[10] [15];
  assign nw02780 = nr00000[1] ? nw02779 : nw02778;
  assign nw02781 = nr00000[0] ? \nr00071[13] [15] : \nr00071[12] [15];
  assign nw02782 = nr00000[0] ? \nr00071[15] [15] : \nr00071[14] [15];
  assign nw02783 = nr00000[1] ? nw02782 : nw02781;
  assign nw02784 = nr00000[2] ? nw02783 : nw02780;
  assign nw02785 = nr00000[3] ? nw02784 : nw02777;
  assign nw02786 = nr00000[0] ? \nr00071[17] [15] : \nr00071[16] [15];
  assign nw02787 = nr00000[0] ? \nr00071[19] [15] : \nr00071[18] [15];
  assign nw02788 = nr00000[1] ? nw02787 : nw02786;
  assign nw02789 = nr00000[0] ? \nr00071[21] [15] : \nr00071[20] [15];
  assign nw02790 = nr00000[0] ? \nr00071[23] [15] : \nr00071[22] [15];
  assign nw02791 = nr00000[1] ? nw02790 : nw02789;
  assign nw02792 = nr00000[2] ? nw02791 : nw02788;
  assign nw02793 = nr00000[0] ? \nr00071[25] [15] : \nr00071[24] [15];
  assign nw02794 = nr00000[0] ? \nr00071[27] [15] : \nr00071[26] [15];
  assign nw02795 = nr00000[1] ? nw02794 : nw02793;
  assign nw02796 = nr00000[0] ? \nr00071[29] [15] : \nr00071[28] [15];
  assign nw02797 = nr00000[0] ? \nr00071[31] [15] : \nr00071[30] [15];
  assign nw02798 = nr00000[1] ? nw02797 : nw02796;
  assign nw02799 = nr00000[2] ? nw02798 : nw02795;
  assign nw02800 = nr00000[3] ? nw02799 : nw02792;
  assign nw00208 = nr00000[4] ? nw02800 : nw02785;
  assign nw02801 = nr00000[0] ? \nr00071[1] [16] : \nr00071[0] [16];
  assign nw02802 = nr00000[0] ? \nr00071[3] [16] : \nr00071[2] [16];
  assign nw02803 = nr00000[1] ? nw02802 : nw02801;
  assign nw02804 = nr00000[0] ? \nr00071[5] [16] : \nr00071[4] [16];
  assign nw02805 = nr00000[0] ? \nr00071[7] [16] : \nr00071[6] [16];
  assign nw02806 = nr00000[1] ? nw02805 : nw02804;
  assign nw02807 = nr00000[2] ? nw02806 : nw02803;
  assign nw02808 = nr00000[0] ? \nr00071[9] [16] : \nr00071[8] [16];
  assign nw02809 = nr00000[0] ? \nr00071[11] [16] : \nr00071[10] [16];
  assign nw02810 = nr00000[1] ? nw02809 : nw02808;
  assign nw02811 = nr00000[0] ? \nr00071[13] [16] : \nr00071[12] [16];
  assign nw02812 = nr00000[0] ? \nr00071[15] [16] : \nr00071[14] [16];
  assign nw02813 = nr00000[1] ? nw02812 : nw02811;
  assign nw02814 = nr00000[2] ? nw02813 : nw02810;
  assign nw02815 = nr00000[3] ? nw02814 : nw02807;
  assign nw02816 = nr00000[0] ? \nr00071[17] [16] : \nr00071[16] [16];
  assign nw02817 = nr00000[0] ? \nr00071[19] [16] : \nr00071[18] [16];
  assign nw02818 = nr00000[1] ? nw02817 : nw02816;
  assign nw02819 = nr00000[0] ? \nr00071[21] [16] : \nr00071[20] [16];
  assign nw02820 = nr00000[0] ? \nr00071[23] [16] : \nr00071[22] [16];
  assign nw02821 = nr00000[1] ? nw02820 : nw02819;
  assign nw02822 = nr00000[2] ? nw02821 : nw02818;
  assign nw02823 = nr00000[0] ? \nr00071[25] [16] : \nr00071[24] [16];
  assign nw02824 = nr00000[0] ? \nr00071[27] [16] : \nr00071[26] [16];
  assign nw02825 = nr00000[1] ? nw02824 : nw02823;
  assign nw02826 = nr00000[0] ? \nr00071[29] [16] : \nr00071[28] [16];
  assign nw02827 = nr00000[0] ? \nr00071[31] [16] : \nr00071[30] [16];
  assign nw02828 = nr00000[1] ? nw02827 : nw02826;
  assign nw02829 = nr00000[2] ? nw02828 : nw02825;
  assign nw02830 = nr00000[3] ? nw02829 : nw02822;
  assign nw00209 = nr00000[4] ? nw02830 : nw02815;
  assign nw02831 = nr00000[0] ? \nr00071[1] [17] : \nr00071[0] [17];
  assign nw02832 = nr00000[0] ? \nr00071[3] [17] : \nr00071[2] [17];
  assign nw02833 = nr00000[1] ? nw02832 : nw02831;
  assign nw02834 = nr00000[0] ? \nr00071[5] [17] : \nr00071[4] [17];
  assign nw02835 = nr00000[0] ? \nr00071[7] [17] : \nr00071[6] [17];
  assign nw02836 = nr00000[1] ? nw02835 : nw02834;
  assign nw02837 = nr00000[2] ? nw02836 : nw02833;
  assign nw02838 = nr00000[0] ? \nr00071[9] [17] : \nr00071[8] [17];
  assign nw02839 = nr00000[0] ? \nr00071[11] [17] : \nr00071[10] [17];
  assign nw02840 = nr00000[1] ? nw02839 : nw02838;
  assign nw02841 = nr00000[0] ? \nr00071[13] [17] : \nr00071[12] [17];
  assign nw02842 = nr00000[0] ? \nr00071[15] [17] : \nr00071[14] [17];
  assign nw02843 = nr00000[1] ? nw02842 : nw02841;
  assign nw02844 = nr00000[2] ? nw02843 : nw02840;
  assign nw02845 = nr00000[3] ? nw02844 : nw02837;
  assign nw02846 = nr00000[0] ? \nr00071[17] [17] : \nr00071[16] [17];
  assign nw02847 = nr00000[0] ? \nr00071[19] [17] : \nr00071[18] [17];
  assign nw02848 = nr00000[1] ? nw02847 : nw02846;
  assign nw02849 = nr00000[0] ? \nr00071[21] [17] : \nr00071[20] [17];
  assign nw02850 = nr00000[0] ? \nr00071[23] [17] : \nr00071[22] [17];
  assign nw02851 = nr00000[1] ? nw02850 : nw02849;
  assign nw02852 = nr00000[2] ? nw02851 : nw02848;
  assign nw02853 = nr00000[0] ? \nr00071[25] [17] : \nr00071[24] [17];
  assign nw02854 = nr00000[0] ? \nr00071[27] [17] : \nr00071[26] [17];
  assign nw02855 = nr00000[1] ? nw02854 : nw02853;
  assign nw02856 = nr00000[0] ? \nr00071[29] [17] : \nr00071[28] [17];
  assign nw02857 = nr00000[0] ? \nr00071[31] [17] : \nr00071[30] [17];
  assign nw02858 = nr00000[1] ? nw02857 : nw02856;
  assign nw02859 = nr00000[2] ? nw02858 : nw02855;
  assign nw02860 = nr00000[3] ? nw02859 : nw02852;
  assign nw00210 = nr00000[4] ? nw02860 : nw02845;
  assign nw02861 = nr00000[0] ? \nr00071[1] [18] : \nr00071[0] [18];
  assign nw02862 = nr00000[0] ? \nr00071[3] [18] : \nr00071[2] [18];
  assign nw02863 = nr00000[1] ? nw02862 : nw02861;
  assign nw02864 = nr00000[0] ? \nr00071[5] [18] : \nr00071[4] [18];
  assign nw02865 = nr00000[0] ? \nr00071[7] [18] : \nr00071[6] [18];
  assign nw02866 = nr00000[1] ? nw02865 : nw02864;
  assign nw02867 = nr00000[2] ? nw02866 : nw02863;
  assign nw02868 = nr00000[0] ? \nr00071[9] [18] : \nr00071[8] [18];
  assign nw02869 = nr00000[0] ? \nr00071[11] [18] : \nr00071[10] [18];
  assign nw02870 = nr00000[1] ? nw02869 : nw02868;
  assign nw02871 = nr00000[0] ? \nr00071[13] [18] : \nr00071[12] [18];
  assign nw02872 = nr00000[0] ? \nr00071[15] [18] : \nr00071[14] [18];
  assign nw02873 = nr00000[1] ? nw02872 : nw02871;
  assign nw02874 = nr00000[2] ? nw02873 : nw02870;
  assign nw02875 = nr00000[3] ? nw02874 : nw02867;
  assign nw02876 = nr00000[0] ? \nr00071[17] [18] : \nr00071[16] [18];
  assign nw02877 = nr00000[0] ? \nr00071[19] [18] : \nr00071[18] [18];
  assign nw02878 = nr00000[1] ? nw02877 : nw02876;
  assign nw02879 = nr00000[0] ? \nr00071[21] [18] : \nr00071[20] [18];
  assign nw02880 = nr00000[0] ? \nr00071[23] [18] : \nr00071[22] [18];
  assign nw02881 = nr00000[1] ? nw02880 : nw02879;
  assign nw02882 = nr00000[2] ? nw02881 : nw02878;
  assign nw02883 = nr00000[0] ? \nr00071[25] [18] : \nr00071[24] [18];
  assign nw02884 = nr00000[0] ? \nr00071[27] [18] : \nr00071[26] [18];
  assign nw02885 = nr00000[1] ? nw02884 : nw02883;
  assign nw02886 = nr00000[0] ? \nr00071[29] [18] : \nr00071[28] [18];
  assign nw02887 = nr00000[0] ? \nr00071[31] [18] : \nr00071[30] [18];
  assign nw02888 = nr00000[1] ? nw02887 : nw02886;
  assign nw02889 = nr00000[2] ? nw02888 : nw02885;
  assign nw02890 = nr00000[3] ? nw02889 : nw02882;
  assign nw00211 = nr00000[4] ? nw02890 : nw02875;
  assign nw02891 = nr00000[0] ? \nr00071[1] [19] : \nr00071[0] [19];
  assign nw02892 = nr00000[0] ? \nr00071[3] [19] : \nr00071[2] [19];
  assign nw02893 = nr00000[1] ? nw02892 : nw02891;
  assign nw02894 = nr00000[0] ? \nr00071[5] [19] : \nr00071[4] [19];
  assign nw02895 = nr00000[0] ? \nr00071[7] [19] : \nr00071[6] [19];
  assign nw02896 = nr00000[1] ? nw02895 : nw02894;
  assign nw02897 = nr00000[2] ? nw02896 : nw02893;
  assign nw02898 = nr00000[0] ? \nr00071[9] [19] : \nr00071[8] [19];
  assign nw02899 = nr00000[0] ? \nr00071[11] [19] : \nr00071[10] [19];
  assign nw02900 = nr00000[1] ? nw02899 : nw02898;
  assign nw02901 = nr00000[0] ? \nr00071[13] [19] : \nr00071[12] [19];
  assign nw02902 = nr00000[0] ? \nr00071[15] [19] : \nr00071[14] [19];
  assign nw02903 = nr00000[1] ? nw02902 : nw02901;
  assign nw02904 = nr00000[2] ? nw02903 : nw02900;
  assign nw02905 = nr00000[3] ? nw02904 : nw02897;
  assign nw02906 = nr00000[0] ? \nr00071[17] [19] : \nr00071[16] [19];
  assign nw02907 = nr00000[0] ? \nr00071[19] [19] : \nr00071[18] [19];
  assign nw02908 = nr00000[1] ? nw02907 : nw02906;
  assign nw02909 = nr00000[0] ? \nr00071[21] [19] : \nr00071[20] [19];
  assign nw02910 = nr00000[0] ? \nr00071[23] [19] : \nr00071[22] [19];
  assign nw02911 = nr00000[1] ? nw02910 : nw02909;
  assign nw02912 = nr00000[2] ? nw02911 : nw02908;
  assign nw02913 = nr00000[0] ? \nr00071[25] [19] : \nr00071[24] [19];
  assign nw02914 = nr00000[0] ? \nr00071[27] [19] : \nr00071[26] [19];
  assign nw02915 = nr00000[1] ? nw02914 : nw02913;
  assign nw02916 = nr00000[0] ? \nr00071[29] [19] : \nr00071[28] [19];
  assign nw02917 = nr00000[0] ? \nr00071[31] [19] : \nr00071[30] [19];
  assign nw02918 = nr00000[1] ? nw02917 : nw02916;
  assign nw02919 = nr00000[2] ? nw02918 : nw02915;
  assign nw02920 = nr00000[3] ? nw02919 : nw02912;
  assign nw00212 = nr00000[4] ? nw02920 : nw02905;
  assign nw02921 = nr00000[0] ? \nr00071[1] [20] : \nr00071[0] [20];
  assign nw02922 = nr00000[0] ? \nr00071[3] [20] : \nr00071[2] [20];
  assign nw02923 = nr00000[1] ? nw02922 : nw02921;
  assign nw02924 = nr00000[0] ? \nr00071[5] [20] : \nr00071[4] [20];
  assign nw02925 = nr00000[0] ? \nr00071[7] [20] : \nr00071[6] [20];
  assign nw02926 = nr00000[1] ? nw02925 : nw02924;
  assign nw02927 = nr00000[2] ? nw02926 : nw02923;
  assign nw02928 = nr00000[0] ? \nr00071[9] [20] : \nr00071[8] [20];
  assign nw02929 = nr00000[0] ? \nr00071[11] [20] : \nr00071[10] [20];
  assign nw02930 = nr00000[1] ? nw02929 : nw02928;
  assign nw02931 = nr00000[0] ? \nr00071[13] [20] : \nr00071[12] [20];
  assign nw02932 = nr00000[0] ? \nr00071[15] [20] : \nr00071[14] [20];
  assign nw02933 = nr00000[1] ? nw02932 : nw02931;
  assign nw02934 = nr00000[2] ? nw02933 : nw02930;
  assign nw02935 = nr00000[3] ? nw02934 : nw02927;
  assign nw02936 = nr00000[0] ? \nr00071[17] [20] : \nr00071[16] [20];
  assign nw02937 = nr00000[0] ? \nr00071[19] [20] : \nr00071[18] [20];
  assign nw02938 = nr00000[1] ? nw02937 : nw02936;
  assign nw02939 = nr00000[0] ? \nr00071[21] [20] : \nr00071[20] [20];
  assign nw02940 = nr00000[0] ? \nr00071[23] [20] : \nr00071[22] [20];
  assign nw02941 = nr00000[1] ? nw02940 : nw02939;
  assign nw02942 = nr00000[2] ? nw02941 : nw02938;
  assign nw02943 = nr00000[0] ? \nr00071[25] [20] : \nr00071[24] [20];
  assign nw02944 = nr00000[0] ? \nr00071[27] [20] : \nr00071[26] [20];
  assign nw02945 = nr00000[1] ? nw02944 : nw02943;
  assign nw02946 = nr00000[0] ? \nr00071[29] [20] : \nr00071[28] [20];
  assign nw02947 = nr00000[0] ? \nr00071[31] [20] : \nr00071[30] [20];
  assign nw02948 = nr00000[1] ? nw02947 : nw02946;
  assign nw02949 = nr00000[2] ? nw02948 : nw02945;
  assign nw02950 = nr00000[3] ? nw02949 : nw02942;
  assign nw00214 = nr00000[4] ? nw02950 : nw02935;
  assign nw02951 = nr00000[0] ? \nr00071[1] [21] : \nr00071[0] [21];
  assign nw02952 = nr00000[0] ? \nr00071[3] [21] : \nr00071[2] [21];
  assign nw02953 = nr00000[1] ? nw02952 : nw02951;
  assign nw02954 = nr00000[0] ? \nr00071[5] [21] : \nr00071[4] [21];
  assign nw02955 = nr00000[0] ? \nr00071[7] [21] : \nr00071[6] [21];
  assign nw02956 = nr00000[1] ? nw02955 : nw02954;
  assign nw02957 = nr00000[2] ? nw02956 : nw02953;
  assign nw02958 = nr00000[0] ? \nr00071[9] [21] : \nr00071[8] [21];
  assign nw02959 = nr00000[0] ? \nr00071[11] [21] : \nr00071[10] [21];
  assign nw02960 = nr00000[1] ? nw02959 : nw02958;
  assign nw02961 = nr00000[0] ? \nr00071[13] [21] : \nr00071[12] [21];
  assign nw02962 = nr00000[0] ? \nr00071[15] [21] : \nr00071[14] [21];
  assign nw02963 = nr00000[1] ? nw02962 : nw02961;
  assign nw02964 = nr00000[2] ? nw02963 : nw02960;
  assign nw02965 = nr00000[3] ? nw02964 : nw02957;
  assign nw02966 = nr00000[0] ? \nr00071[17] [21] : \nr00071[16] [21];
  assign nw02967 = nr00000[0] ? \nr00071[19] [21] : \nr00071[18] [21];
  assign nw02968 = nr00000[1] ? nw02967 : nw02966;
  assign nw02969 = nr00000[0] ? \nr00071[21] [21] : \nr00071[20] [21];
  assign nw02970 = nr00000[0] ? \nr00071[23] [21] : \nr00071[22] [21];
  assign nw02971 = nr00000[1] ? nw02970 : nw02969;
  assign nw02972 = nr00000[2] ? nw02971 : nw02968;
  assign nw02973 = nr00000[0] ? \nr00071[25] [21] : \nr00071[24] [21];
  assign nw02974 = nr00000[0] ? \nr00071[27] [21] : \nr00071[26] [21];
  assign nw02975 = nr00000[1] ? nw02974 : nw02973;
  assign nw02976 = nr00000[0] ? \nr00071[29] [21] : \nr00071[28] [21];
  assign nw02977 = nr00000[0] ? \nr00071[31] [21] : \nr00071[30] [21];
  assign nw02978 = nr00000[1] ? nw02977 : nw02976;
  assign nw02979 = nr00000[2] ? nw02978 : nw02975;
  assign nw02980 = nr00000[3] ? nw02979 : nw02972;
  assign nw00215 = nr00000[4] ? nw02980 : nw02965;
  assign nw02981 = nr00000[0] ? \nr00071[1] [22] : \nr00071[0] [22];
  assign nw02982 = nr00000[0] ? \nr00071[3] [22] : \nr00071[2] [22];
  assign nw02983 = nr00000[1] ? nw02982 : nw02981;
  assign nw02984 = nr00000[0] ? \nr00071[5] [22] : \nr00071[4] [22];
  assign nw02985 = nr00000[0] ? \nr00071[7] [22] : \nr00071[6] [22];
  assign nw02986 = nr00000[1] ? nw02985 : nw02984;
  assign nw02987 = nr00000[2] ? nw02986 : nw02983;
  assign nw02988 = nr00000[0] ? \nr00071[9] [22] : \nr00071[8] [22];
  assign nw02989 = nr00000[0] ? \nr00071[11] [22] : \nr00071[10] [22];
  assign nw02990 = nr00000[1] ? nw02989 : nw02988;
  assign nw02991 = nr00000[0] ? \nr00071[13] [22] : \nr00071[12] [22];
  assign nw02992 = nr00000[0] ? \nr00071[15] [22] : \nr00071[14] [22];
  assign nw02993 = nr00000[1] ? nw02992 : nw02991;
  assign nw02994 = nr00000[2] ? nw02993 : nw02990;
  assign nw02995 = nr00000[3] ? nw02994 : nw02987;
  assign nw02996 = nr00000[0] ? \nr00071[17] [22] : \nr00071[16] [22];
  assign nw02997 = nr00000[0] ? \nr00071[19] [22] : \nr00071[18] [22];
  assign nw02998 = nr00000[1] ? nw02997 : nw02996;
  assign nw02999 = nr00000[0] ? \nr00071[21] [22] : \nr00071[20] [22];
  assign nw03000 = nr00000[0] ? \nr00071[23] [22] : \nr00071[22] [22];
  assign nw03001 = nr00000[1] ? nw03000 : nw02999;
  assign nw03002 = nr00000[2] ? nw03001 : nw02998;
  assign nw03003 = nr00000[0] ? \nr00071[25] [22] : \nr00071[24] [22];
  assign nw03004 = nr00000[0] ? \nr00071[27] [22] : \nr00071[26] [22];
  assign nw03005 = nr00000[1] ? nw03004 : nw03003;
  assign nw03006 = nr00000[0] ? \nr00071[29] [22] : \nr00071[28] [22];
  assign nw03007 = nr00000[0] ? \nr00071[31] [22] : \nr00071[30] [22];
  assign nw03008 = nr00000[1] ? nw03007 : nw03006;
  assign nw03009 = nr00000[2] ? nw03008 : nw03005;
  assign nw03010 = nr00000[3] ? nw03009 : nw03002;
  assign nw00216 = nr00000[4] ? nw03010 : nw02995;
  assign nw03011 = nr00000[0] ? \nr00071[1] [23] : \nr00071[0] [23];
  assign nw03012 = nr00000[0] ? \nr00071[3] [23] : \nr00071[2] [23];
  assign nw03013 = nr00000[1] ? nw03012 : nw03011;
  assign nw03014 = nr00000[0] ? \nr00071[5] [23] : \nr00071[4] [23];
  assign nw03015 = nr00000[0] ? \nr00071[7] [23] : \nr00071[6] [23];
  assign nw03016 = nr00000[1] ? nw03015 : nw03014;
  assign nw03017 = nr00000[2] ? nw03016 : nw03013;
  assign nw03018 = nr00000[0] ? \nr00071[9] [23] : \nr00071[8] [23];
  assign nw03019 = nr00000[0] ? \nr00071[11] [23] : \nr00071[10] [23];
  assign nw03020 = nr00000[1] ? nw03019 : nw03018;
  assign nw03021 = nr00000[0] ? \nr00071[13] [23] : \nr00071[12] [23];
  assign nw03022 = nr00000[0] ? \nr00071[15] [23] : \nr00071[14] [23];
  assign nw03023 = nr00000[1] ? nw03022 : nw03021;
  assign nw03024 = nr00000[2] ? nw03023 : nw03020;
  assign nw03025 = nr00000[3] ? nw03024 : nw03017;
  assign nw03026 = nr00000[0] ? \nr00071[17] [23] : \nr00071[16] [23];
  assign nw03027 = nr00000[0] ? \nr00071[19] [23] : \nr00071[18] [23];
  assign nw03028 = nr00000[1] ? nw03027 : nw03026;
  assign nw03029 = nr00000[0] ? \nr00071[21] [23] : \nr00071[20] [23];
  assign nw03030 = nr00000[0] ? \nr00071[23] [23] : \nr00071[22] [23];
  assign nw03031 = nr00000[1] ? nw03030 : nw03029;
  assign nw03032 = nr00000[2] ? nw03031 : nw03028;
  assign nw03033 = nr00000[0] ? \nr00071[25] [23] : \nr00071[24] [23];
  assign nw03034 = nr00000[0] ? \nr00071[27] [23] : \nr00071[26] [23];
  assign nw03035 = nr00000[1] ? nw03034 : nw03033;
  assign nw03036 = nr00000[0] ? \nr00071[29] [23] : \nr00071[28] [23];
  assign nw03037 = nr00000[0] ? \nr00071[31] [23] : \nr00071[30] [23];
  assign nw03038 = nr00000[1] ? nw03037 : nw03036;
  assign nw03039 = nr00000[2] ? nw03038 : nw03035;
  assign nw03040 = nr00000[3] ? nw03039 : nw03032;
  assign nw00217 = nr00000[4] ? nw03040 : nw03025;
  assign nw03041 = nr00000[0] ? \nr00071[1] [24] : \nr00071[0] [24];
  assign nw03042 = nr00000[0] ? \nr00071[3] [24] : \nr00071[2] [24];
  assign nw03043 = nr00000[1] ? nw03042 : nw03041;
  assign nw03044 = nr00000[0] ? \nr00071[5] [24] : \nr00071[4] [24];
  assign nw03045 = nr00000[0] ? \nr00071[7] [24] : \nr00071[6] [24];
  assign nw03046 = nr00000[1] ? nw03045 : nw03044;
  assign nw03047 = nr00000[2] ? nw03046 : nw03043;
  assign nw03048 = nr00000[0] ? \nr00071[9] [24] : \nr00071[8] [24];
  assign nw03049 = nr00000[0] ? \nr00071[11] [24] : \nr00071[10] [24];
  assign nw03050 = nr00000[1] ? nw03049 : nw03048;
  assign nw03051 = nr00000[0] ? \nr00071[13] [24] : \nr00071[12] [24];
  assign nw03052 = nr00000[0] ? \nr00071[15] [24] : \nr00071[14] [24];
  assign nw03053 = nr00000[1] ? nw03052 : nw03051;
  assign nw03054 = nr00000[2] ? nw03053 : nw03050;
  assign nw03055 = nr00000[3] ? nw03054 : nw03047;
  assign nw03056 = nr00000[0] ? \nr00071[17] [24] : \nr00071[16] [24];
  assign nw03057 = nr00000[0] ? \nr00071[19] [24] : \nr00071[18] [24];
  assign nw03058 = nr00000[1] ? nw03057 : nw03056;
  assign nw03059 = nr00000[0] ? \nr00071[21] [24] : \nr00071[20] [24];
  assign nw03060 = nr00000[0] ? \nr00071[23] [24] : \nr00071[22] [24];
  assign nw03061 = nr00000[1] ? nw03060 : nw03059;
  assign nw03062 = nr00000[2] ? nw03061 : nw03058;
  assign nw03063 = nr00000[0] ? \nr00071[25] [24] : \nr00071[24] [24];
  assign nw03064 = nr00000[0] ? \nr00071[27] [24] : \nr00071[26] [24];
  assign nw03065 = nr00000[1] ? nw03064 : nw03063;
  assign nw03066 = nr00000[0] ? \nr00071[29] [24] : \nr00071[28] [24];
  assign nw03067 = nr00000[0] ? \nr00071[31] [24] : \nr00071[30] [24];
  assign nw03068 = nr00000[1] ? nw03067 : nw03066;
  assign nw03069 = nr00000[2] ? nw03068 : nw03065;
  assign nw03070 = nr00000[3] ? nw03069 : nw03062;
  assign nw00218 = nr00000[4] ? nw03070 : nw03055;
  assign nw03071 = nr00000[0] ? \nr00071[1] [25] : \nr00071[0] [25];
  assign nw03072 = nr00000[0] ? \nr00071[3] [25] : \nr00071[2] [25];
  assign nw03073 = nr00000[1] ? nw03072 : nw03071;
  assign nw03074 = nr00000[0] ? \nr00071[5] [25] : \nr00071[4] [25];
  assign nw03075 = nr00000[0] ? \nr00071[7] [25] : \nr00071[6] [25];
  assign nw03076 = nr00000[1] ? nw03075 : nw03074;
  assign nw03077 = nr00000[2] ? nw03076 : nw03073;
  assign nw03078 = nr00000[0] ? \nr00071[9] [25] : \nr00071[8] [25];
  assign nw03079 = nr00000[0] ? \nr00071[11] [25] : \nr00071[10] [25];
  assign nw03080 = nr00000[1] ? nw03079 : nw03078;
  assign nw03081 = nr00000[0] ? \nr00071[13] [25] : \nr00071[12] [25];
  assign nw03082 = nr00000[0] ? \nr00071[15] [25] : \nr00071[14] [25];
  assign nw03083 = nr00000[1] ? nw03082 : nw03081;
  assign nw03084 = nr00000[2] ? nw03083 : nw03080;
  assign nw03085 = nr00000[3] ? nw03084 : nw03077;
  assign nw03086 = nr00000[0] ? \nr00071[17] [25] : \nr00071[16] [25];
  assign nw03087 = nr00000[0] ? \nr00071[19] [25] : \nr00071[18] [25];
  assign nw03088 = nr00000[1] ? nw03087 : nw03086;
  assign nw03089 = nr00000[0] ? \nr00071[21] [25] : \nr00071[20] [25];
  assign nw03090 = nr00000[0] ? \nr00071[23] [25] : \nr00071[22] [25];
  assign nw03091 = nr00000[1] ? nw03090 : nw03089;
  assign nw03092 = nr00000[2] ? nw03091 : nw03088;
  assign nw03093 = nr00000[0] ? \nr00071[25] [25] : \nr00071[24] [25];
  assign nw03094 = nr00000[0] ? \nr00071[27] [25] : \nr00071[26] [25];
  assign nw03095 = nr00000[1] ? nw03094 : nw03093;
  assign nw03096 = nr00000[0] ? \nr00071[29] [25] : \nr00071[28] [25];
  assign nw03097 = nr00000[0] ? \nr00071[31] [25] : \nr00071[30] [25];
  assign nw03098 = nr00000[1] ? nw03097 : nw03096;
  assign nw03099 = nr00000[2] ? nw03098 : nw03095;
  assign nw03100 = nr00000[3] ? nw03099 : nw03092;
  assign nw00219 = nr00000[4] ? nw03100 : nw03085;
  assign nw03101 = nr00000[0] ? \nr00071[1] [26] : \nr00071[0] [26];
  assign nw03102 = nr00000[0] ? \nr00071[3] [26] : \nr00071[2] [26];
  assign nw03103 = nr00000[1] ? nw03102 : nw03101;
  assign nw03104 = nr00000[0] ? \nr00071[5] [26] : \nr00071[4] [26];
  assign nw03105 = nr00000[0] ? \nr00071[7] [26] : \nr00071[6] [26];
  assign nw03106 = nr00000[1] ? nw03105 : nw03104;
  assign nw03107 = nr00000[2] ? nw03106 : nw03103;
  assign nw03108 = nr00000[0] ? \nr00071[9] [26] : \nr00071[8] [26];
  assign nw03109 = nr00000[0] ? \nr00071[11] [26] : \nr00071[10] [26];
  assign nw03110 = nr00000[1] ? nw03109 : nw03108;
  assign nw03111 = nr00000[0] ? \nr00071[13] [26] : \nr00071[12] [26];
  assign nw03112 = nr00000[0] ? \nr00071[15] [26] : \nr00071[14] [26];
  assign nw03113 = nr00000[1] ? nw03112 : nw03111;
  assign nw03114 = nr00000[2] ? nw03113 : nw03110;
  assign nw03115 = nr00000[3] ? nw03114 : nw03107;
  assign nw03116 = nr00000[0] ? \nr00071[17] [26] : \nr00071[16] [26];
  assign nw03117 = nr00000[0] ? \nr00071[19] [26] : \nr00071[18] [26];
  assign nw03118 = nr00000[1] ? nw03117 : nw03116;
  assign nw03119 = nr00000[0] ? \nr00071[21] [26] : \nr00071[20] [26];
  assign nw03120 = nr00000[0] ? \nr00071[23] [26] : \nr00071[22] [26];
  assign nw03121 = nr00000[1] ? nw03120 : nw03119;
  assign nw03122 = nr00000[2] ? nw03121 : nw03118;
  assign nw03123 = nr00000[0] ? \nr00071[25] [26] : \nr00071[24] [26];
  assign nw03124 = nr00000[0] ? \nr00071[27] [26] : \nr00071[26] [26];
  assign nw03125 = nr00000[1] ? nw03124 : nw03123;
  assign nw03126 = nr00000[0] ? \nr00071[29] [26] : \nr00071[28] [26];
  assign nw03127 = nr00000[0] ? \nr00071[31] [26] : \nr00071[30] [26];
  assign nw03128 = nr00000[1] ? nw03127 : nw03126;
  assign nw03129 = nr00000[2] ? nw03128 : nw03125;
  assign nw03130 = nr00000[3] ? nw03129 : nw03122;
  assign nw00220 = nr00000[4] ? nw03130 : nw03115;
  assign nw03131 = nr00000[0] ? \nr00071[1] [27] : \nr00071[0] [27];
  assign nw03132 = nr00000[0] ? \nr00071[3] [27] : \nr00071[2] [27];
  assign nw03133 = nr00000[1] ? nw03132 : nw03131;
  assign nw03134 = nr00000[0] ? \nr00071[5] [27] : \nr00071[4] [27];
  assign nw03135 = nr00000[0] ? \nr00071[7] [27] : \nr00071[6] [27];
  assign nw03136 = nr00000[1] ? nw03135 : nw03134;
  assign nw03137 = nr00000[2] ? nw03136 : nw03133;
  assign nw03138 = nr00000[0] ? \nr00071[9] [27] : \nr00071[8] [27];
  assign nw03139 = nr00000[0] ? \nr00071[11] [27] : \nr00071[10] [27];
  assign nw03140 = nr00000[1] ? nw03139 : nw03138;
  assign nw03141 = nr00000[0] ? \nr00071[13] [27] : \nr00071[12] [27];
  assign nw03142 = nr00000[0] ? \nr00071[15] [27] : \nr00071[14] [27];
  assign nw03143 = nr00000[1] ? nw03142 : nw03141;
  assign nw03144 = nr00000[2] ? nw03143 : nw03140;
  assign nw03145 = nr00000[3] ? nw03144 : nw03137;
  assign nw03146 = nr00000[0] ? \nr00071[17] [27] : \nr00071[16] [27];
  assign nw03147 = nr00000[0] ? \nr00071[19] [27] : \nr00071[18] [27];
  assign nw03148 = nr00000[1] ? nw03147 : nw03146;
  assign nw03149 = nr00000[0] ? \nr00071[21] [27] : \nr00071[20] [27];
  assign nw03150 = nr00000[0] ? \nr00071[23] [27] : \nr00071[22] [27];
  assign nw03151 = nr00000[1] ? nw03150 : nw03149;
  assign nw03152 = nr00000[2] ? nw03151 : nw03148;
  assign nw03153 = nr00000[0] ? \nr00071[25] [27] : \nr00071[24] [27];
  assign nw03154 = nr00000[0] ? \nr00071[27] [27] : \nr00071[26] [27];
  assign nw03155 = nr00000[1] ? nw03154 : nw03153;
  assign nw03156 = nr00000[0] ? \nr00071[29] [27] : \nr00071[28] [27];
  assign nw03157 = nr00000[0] ? \nr00071[31] [27] : \nr00071[30] [27];
  assign nw03158 = nr00000[1] ? nw03157 : nw03156;
  assign nw03159 = nr00000[2] ? nw03158 : nw03155;
  assign nw03160 = nr00000[3] ? nw03159 : nw03152;
  assign nw00221 = nr00000[4] ? nw03160 : nw03145;
  assign nw03161 = nr00000[0] ? \nr00071[1] [28] : \nr00071[0] [28];
  assign nw03162 = nr00000[0] ? \nr00071[3] [28] : \nr00071[2] [28];
  assign nw03163 = nr00000[1] ? nw03162 : nw03161;
  assign nw03164 = nr00000[0] ? \nr00071[5] [28] : \nr00071[4] [28];
  assign nw03165 = nr00000[0] ? \nr00071[7] [28] : \nr00071[6] [28];
  assign nw03166 = nr00000[1] ? nw03165 : nw03164;
  assign nw03167 = nr00000[2] ? nw03166 : nw03163;
  assign nw03168 = nr00000[0] ? \nr00071[9] [28] : \nr00071[8] [28];
  assign nw03169 = nr00000[0] ? \nr00071[11] [28] : \nr00071[10] [28];
  assign nw03170 = nr00000[1] ? nw03169 : nw03168;
  assign nw03171 = nr00000[0] ? \nr00071[13] [28] : \nr00071[12] [28];
  assign nw03172 = nr00000[0] ? \nr00071[15] [28] : \nr00071[14] [28];
  assign nw03173 = nr00000[1] ? nw03172 : nw03171;
  assign nw03174 = nr00000[2] ? nw03173 : nw03170;
  assign nw03175 = nr00000[3] ? nw03174 : nw03167;
  assign nw03176 = nr00000[0] ? \nr00071[17] [28] : \nr00071[16] [28];
  assign nw03177 = nr00000[0] ? \nr00071[19] [28] : \nr00071[18] [28];
  assign nw03178 = nr00000[1] ? nw03177 : nw03176;
  assign nw03179 = nr00000[0] ? \nr00071[21] [28] : \nr00071[20] [28];
  assign nw03180 = nr00000[0] ? \nr00071[23] [28] : \nr00071[22] [28];
  assign nw03181 = nr00000[1] ? nw03180 : nw03179;
  assign nw03182 = nr00000[2] ? nw03181 : nw03178;
  assign nw03183 = nr00000[0] ? \nr00071[25] [28] : \nr00071[24] [28];
  assign nw03184 = nr00000[0] ? \nr00071[27] [28] : \nr00071[26] [28];
  assign nw03185 = nr00000[1] ? nw03184 : nw03183;
  assign nw03186 = nr00000[0] ? \nr00071[29] [28] : \nr00071[28] [28];
  assign nw03187 = nr00000[0] ? \nr00071[31] [28] : \nr00071[30] [28];
  assign nw03188 = nr00000[1] ? nw03187 : nw03186;
  assign nw03189 = nr00000[2] ? nw03188 : nw03185;
  assign nw03190 = nr00000[3] ? nw03189 : nw03182;
  assign nw00222 = nr00000[4] ? nw03190 : nw03175;
  assign nw03191 = nr00000[0] ? \nr00071[1] [29] : \nr00071[0] [29];
  assign nw03192 = nr00000[0] ? \nr00071[3] [29] : \nr00071[2] [29];
  assign nw03193 = nr00000[1] ? nw03192 : nw03191;
  assign nw03194 = nr00000[0] ? \nr00071[5] [29] : \nr00071[4] [29];
  assign nw03195 = nr00000[0] ? \nr00071[7] [29] : \nr00071[6] [29];
  assign nw03196 = nr00000[1] ? nw03195 : nw03194;
  assign nw03197 = nr00000[2] ? nw03196 : nw03193;
  assign nw03198 = nr00000[0] ? \nr00071[9] [29] : \nr00071[8] [29];
  assign nw03199 = nr00000[0] ? \nr00071[11] [29] : \nr00071[10] [29];
  assign nw03200 = nr00000[1] ? nw03199 : nw03198;
  assign nw03201 = nr00000[0] ? \nr00071[13] [29] : \nr00071[12] [29];
  assign nw03202 = nr00000[0] ? \nr00071[15] [29] : \nr00071[14] [29];
  assign nw03203 = nr00000[1] ? nw03202 : nw03201;
  assign nw03204 = nr00000[2] ? nw03203 : nw03200;
  assign nw03205 = nr00000[3] ? nw03204 : nw03197;
  assign nw03206 = nr00000[0] ? \nr00071[17] [29] : \nr00071[16] [29];
  assign nw03207 = nr00000[0] ? \nr00071[19] [29] : \nr00071[18] [29];
  assign nw03208 = nr00000[1] ? nw03207 : nw03206;
  assign nw03209 = nr00000[0] ? \nr00071[21] [29] : \nr00071[20] [29];
  assign nw03210 = nr00000[0] ? \nr00071[23] [29] : \nr00071[22] [29];
  assign nw03211 = nr00000[1] ? nw03210 : nw03209;
  assign nw03212 = nr00000[2] ? nw03211 : nw03208;
  assign nw03213 = nr00000[0] ? \nr00071[25] [29] : \nr00071[24] [29];
  assign nw03214 = nr00000[0] ? \nr00071[27] [29] : \nr00071[26] [29];
  assign nw03215 = nr00000[1] ? nw03214 : nw03213;
  assign nw03216 = nr00000[0] ? \nr00071[29] [29] : \nr00071[28] [29];
  assign nw03217 = nr00000[0] ? \nr00071[31] [29] : \nr00071[30] [29];
  assign nw03218 = nr00000[1] ? nw03217 : nw03216;
  assign nw03219 = nr00000[2] ? nw03218 : nw03215;
  assign nw03220 = nr00000[3] ? nw03219 : nw03212;
  assign nw00223 = nr00000[4] ? nw03220 : nw03205;
  assign nw03221 = nr00000[0] ? \nr00071[1] [30] : \nr00071[0] [30];
  assign nw03222 = nr00000[0] ? \nr00071[3] [30] : \nr00071[2] [30];
  assign nw03223 = nr00000[1] ? nw03222 : nw03221;
  assign nw03224 = nr00000[0] ? \nr00071[5] [30] : \nr00071[4] [30];
  assign nw03225 = nr00000[0] ? \nr00071[7] [30] : \nr00071[6] [30];
  assign nw03226 = nr00000[1] ? nw03225 : nw03224;
  assign nw03227 = nr00000[2] ? nw03226 : nw03223;
  assign nw03228 = nr00000[0] ? \nr00071[9] [30] : \nr00071[8] [30];
  assign nw03229 = nr00000[0] ? \nr00071[11] [30] : \nr00071[10] [30];
  assign nw03230 = nr00000[1] ? nw03229 : nw03228;
  assign nw03231 = nr00000[0] ? \nr00071[13] [30] : \nr00071[12] [30];
  assign nw03232 = nr00000[0] ? \nr00071[15] [30] : \nr00071[14] [30];
  assign nw03233 = nr00000[1] ? nw03232 : nw03231;
  assign nw03234 = nr00000[2] ? nw03233 : nw03230;
  assign nw03235 = nr00000[3] ? nw03234 : nw03227;
  assign nw03236 = nr00000[0] ? \nr00071[17] [30] : \nr00071[16] [30];
  assign nw03237 = nr00000[0] ? \nr00071[19] [30] : \nr00071[18] [30];
  assign nw03238 = nr00000[1] ? nw03237 : nw03236;
  assign nw03239 = nr00000[0] ? \nr00071[21] [30] : \nr00071[20] [30];
  assign nw03240 = nr00000[0] ? \nr00071[23] [30] : \nr00071[22] [30];
  assign nw03241 = nr00000[1] ? nw03240 : nw03239;
  assign nw03242 = nr00000[2] ? nw03241 : nw03238;
  assign nw03243 = nr00000[0] ? \nr00071[25] [30] : \nr00071[24] [30];
  assign nw03244 = nr00000[0] ? \nr00071[27] [30] : \nr00071[26] [30];
  assign nw03245 = nr00000[1] ? nw03244 : nw03243;
  assign nw03246 = nr00000[0] ? \nr00071[29] [30] : \nr00071[28] [30];
  assign nw03247 = nr00000[0] ? \nr00071[31] [30] : \nr00071[30] [30];
  assign nw03248 = nr00000[1] ? nw03247 : nw03246;
  assign nw03249 = nr00000[2] ? nw03248 : nw03245;
  assign nw03250 = nr00000[3] ? nw03249 : nw03242;
  assign nw00225 = nr00000[4] ? nw03250 : nw03235;
  assign nw03251 = nr00000[0] ? \nr00071[1] [31] : \nr00071[0] [31];
  assign nw03252 = nr00000[0] ? \nr00071[3] [31] : \nr00071[2] [31];
  assign nw03253 = nr00000[1] ? nw03252 : nw03251;
  assign nw03254 = nr00000[0] ? \nr00071[5] [31] : \nr00071[4] [31];
  assign nw03255 = nr00000[0] ? \nr00071[7] [31] : \nr00071[6] [31];
  assign nw03256 = nr00000[1] ? nw03255 : nw03254;
  assign nw03257 = nr00000[2] ? nw03256 : nw03253;
  assign nw03258 = nr00000[0] ? \nr00071[9] [31] : \nr00071[8] [31];
  assign nw03259 = nr00000[0] ? \nr00071[11] [31] : \nr00071[10] [31];
  assign nw03260 = nr00000[1] ? nw03259 : nw03258;
  assign nw03261 = nr00000[0] ? \nr00071[13] [31] : \nr00071[12] [31];
  assign nw03262 = nr00000[0] ? \nr00071[15] [31] : \nr00071[14] [31];
  assign nw03263 = nr00000[1] ? nw03262 : nw03261;
  assign nw03264 = nr00000[2] ? nw03263 : nw03260;
  assign nw03265 = nr00000[3] ? nw03264 : nw03257;
  assign nw03266 = nr00000[0] ? \nr00071[17] [31] : \nr00071[16] [31];
  assign nw03267 = nr00000[0] ? \nr00071[19] [31] : \nr00071[18] [31];
  assign nw03268 = nr00000[1] ? nw03267 : nw03266;
  assign nw03269 = nr00000[0] ? \nr00071[21] [31] : \nr00071[20] [31];
  assign nw03270 = nr00000[0] ? \nr00071[23] [31] : \nr00071[22] [31];
  assign nw03271 = nr00000[1] ? nw03270 : nw03269;
  assign nw03272 = nr00000[2] ? nw03271 : nw03268;
  assign nw03273 = nr00000[0] ? \nr00071[25] [31] : \nr00071[24] [31];
  assign nw03274 = nr00000[0] ? \nr00071[27] [31] : \nr00071[26] [31];
  assign nw03275 = nr00000[1] ? nw03274 : nw03273;
  assign nw03276 = nr00000[0] ? \nr00071[29] [31] : \nr00071[28] [31];
  assign nw03277 = nr00000[0] ? \nr00071[31] [31] : \nr00071[30] [31];
  assign nw03278 = nr00000[1] ? nw03277 : nw03276;
  assign nw03279 = nr00000[2] ? nw03278 : nw03275;
  assign nw03280 = nr00000[3] ? nw03279 : nw03272;
  assign nw00226 = nr00000[4] ? nw03280 : nw03265;
  assign nw03281 = \nr00065  & ~(\nr00063 );
  assign nw03282 = nw03281 | ~(nw00656);
  assign nw00383 = \nr00063  ? nw03281 : nw03282;
  assign nw00351 = \nr00025 [1] ? nw01388 : \nr00066 [0];
  assign nw00362 = \nr00025 [1] ? nw01416 : \nr00066 [1];
  assign nw00373 = \nr00025 [1] ? nw01444 : \nr00066 [2];
  assign nw00376 = \nr00025 [1] ? nw01472 : \nr00066 [3];
  assign nw00377 = \nr00025 [1] ? nw01500 : \nr00066 [4];
  assign nw00378 = \nr00025 [1] ? nw01528 : \nr00066 [5];
  assign nw00379 = \nr00025 [1] ? nw01556 : \nr00066 [6];
  assign nw00380 = \nr00025 [1] ? nw01584 : \nr00066 [7];
  assign nw00381 = \nr00025 [1] ? nw01620 : \nr00066 [8];
  assign nw00382 = \nr00025 [1] ? nw01653 : \nr00066 [9];
  assign nw00352 = \nr00025 [1] ? nw01686 : \nr00066 [10];
  assign nw00353 = \nr00025 [1] ? nw01719 : \nr00066 [11];
  assign nw00354 = \nr00025 [1] ? nw01752 : \nr00066 [12];
  assign nw00355 = \nr00025 [1] ? nw01785 : \nr00066 [13];
  assign nw00356 = \nr00025 [1] ? nw01818 : \nr00066 [14];
  assign nw00357 = \nr00025 [1] ? nw01849 : \nr00066 [15];
  assign nw00358 = \nr00025 [1] ? nw01879 : \nr00066 [16];
  assign nw00359 = \nr00025 [1] ? nw01909 : \nr00066 [17];
  assign nw00360 = \nr00025 [1] ? nw01939 : \nr00066 [18];
  assign nw00361 = \nr00025 [1] ? nw01969 : \nr00066 [19];
  assign nw00363 = \nr00025 [1] ? nw01999 : \nr00066 [20];
  assign nw00364 = \nr00025 [1] ? nw02029 : \nr00066 [21];
  assign nw00365 = \nr00025 [1] ? nw02059 : \nr00066 [22];
  assign nw00366 = \nr00025 [1] ? nw02088 : \nr00066 [23];
  assign nw00367 = \nr00025 [1] ? nw02117 : \nr00066 [24];
  assign nw00368 = \nr00025 [1] ? nw02146 : \nr00066 [25];
  assign nw00369 = \nr00025 [1] ? nw02175 : \nr00066 [26];
  assign nw00370 = \nr00025 [1] ? nw02204 : \nr00066 [27];
  assign nw00371 = \nr00025 [1] ? nw02233 : \nr00066 [28];
  assign nw00372 = \nr00025 [1] ? nw02262 : \nr00066 [29];
  assign nw00374 = \nr00025 [1] ? nw02291 : \nr00066 [30];
  assign nw00375 = \nr00025 [1] ? nw02320 : \nr00066 [31];
  assign nw03283 = nr00008 & ~(nw00657);
  assign nw03284 = ~nw01416;
  assign nw03285 = ~(nw01416 | nw01388);
  assign nw03286 = \nr00048  ? nw03285 : nw03283;
  assign nw03287 = \nr00049  ? nw03284 : nw03286;
  assign nw03288 = nw03287 | \nr00060 ;
  assign nw03289 = \nr00025 [1] ? nw03288 : nw03283;
  assign nw00350 = \nr00063  ? nw03283 : nw03289;
  assign nw03290 = ~\nr00065 ;
  assign nw03291 = ~nw00656;
  assign nw00349 = \nr00063  ? nw03290 : nw03291;
  assign nw03292 = nr00001[0] ? \nr00071[1] [0] : \nr00071[0] [0];
  assign nw03293 = nr00001[0] ? \nr00071[3] [0] : \nr00071[2] [0];
  assign nw03294 = nr00001[1] ? nw03293 : nw03292;
  assign nw03295 = nr00001[0] ? \nr00071[5] [0] : \nr00071[4] [0];
  assign nw03296 = nr00001[0] ? \nr00071[7] [0] : \nr00071[6] [0];
  assign nw03297 = nr00001[1] ? nw03296 : nw03295;
  assign nw03298 = nr00001[2] ? nw03297 : nw03294;
  assign nw03299 = nr00001[0] ? \nr00071[9] [0] : \nr00071[8] [0];
  assign nw03300 = nr00001[0] ? \nr00071[11] [0] : \nr00071[10] [0];
  assign nw03301 = nr00001[1] ? nw03300 : nw03299;
  assign nw03302 = nr00001[0] ? \nr00071[13] [0] : \nr00071[12] [0];
  assign nw03303 = nr00001[0] ? \nr00071[15] [0] : \nr00071[14] [0];
  assign nw03304 = nr00001[1] ? nw03303 : nw03302;
  assign nw03305 = nr00001[2] ? nw03304 : nw03301;
  assign nw03306 = nr00001[3] ? nw03305 : nw03298;
  assign nw03307 = nr00001[0] ? \nr00071[17] [0] : \nr00071[16] [0];
  assign nw03308 = nr00001[0] ? \nr00071[19] [0] : \nr00071[18] [0];
  assign nw03309 = nr00001[1] ? nw03308 : nw03307;
  assign nw03310 = nr00001[0] ? \nr00071[21] [0] : \nr00071[20] [0];
  assign nw03311 = nr00001[0] ? \nr00071[23] [0] : \nr00071[22] [0];
  assign nw03312 = nr00001[1] ? nw03311 : nw03310;
  assign nw03313 = nr00001[2] ? nw03312 : nw03309;
  assign nw03314 = nr00001[0] ? \nr00071[25] [0] : \nr00071[24] [0];
  assign nw03315 = nr00001[0] ? \nr00071[27] [0] : \nr00071[26] [0];
  assign nw03316 = nr00001[1] ? nw03315 : nw03314;
  assign nw03317 = nr00001[0] ? \nr00071[29] [0] : \nr00071[28] [0];
  assign nw03318 = nr00001[0] ? \nr00071[31] [0] : \nr00071[30] [0];
  assign nw03319 = nr00001[1] ? nw03318 : nw03317;
  assign nw03320 = nr00001[2] ? nw03319 : nw03316;
  assign nw03321 = nr00001[3] ? nw03320 : nw03313;
  assign nw00170 = nr00001[4] ? nw03321 : nw03306;
  assign nw03322 = \nr00030  | \nr00038 ;
  assign nw03323 = nw03322 | nw00460;
  assign nw00317 = nw03323 ? \nr00067 [0] : nw00170;
  assign nw03324 = nr00001[0] ? \nr00071[1] [1] : \nr00071[0] [1];
  assign nw03325 = nr00001[0] ? \nr00071[3] [1] : \nr00071[2] [1];
  assign nw03326 = nr00001[1] ? nw03325 : nw03324;
  assign nw03327 = nr00001[0] ? \nr00071[5] [1] : \nr00071[4] [1];
  assign nw03328 = nr00001[0] ? \nr00071[7] [1] : \nr00071[6] [1];
  assign nw03329 = nr00001[1] ? nw03328 : nw03327;
  assign nw03330 = nr00001[2] ? nw03329 : nw03326;
  assign nw03331 = nr00001[0] ? \nr00071[9] [1] : \nr00071[8] [1];
  assign nw03332 = nr00001[0] ? \nr00071[11] [1] : \nr00071[10] [1];
  assign nw03333 = nr00001[1] ? nw03332 : nw03331;
  assign nw03334 = nr00001[0] ? \nr00071[13] [1] : \nr00071[12] [1];
  assign nw03335 = nr00001[0] ? \nr00071[15] [1] : \nr00071[14] [1];
  assign nw03336 = nr00001[1] ? nw03335 : nw03334;
  assign nw03337 = nr00001[2] ? nw03336 : nw03333;
  assign nw03338 = nr00001[3] ? nw03337 : nw03330;
  assign nw03339 = nr00001[0] ? \nr00071[17] [1] : \nr00071[16] [1];
  assign nw03340 = nr00001[0] ? \nr00071[19] [1] : \nr00071[18] [1];
  assign nw03341 = nr00001[1] ? nw03340 : nw03339;
  assign nw03342 = nr00001[0] ? \nr00071[21] [1] : \nr00071[20] [1];
  assign nw03343 = nr00001[0] ? \nr00071[23] [1] : \nr00071[22] [1];
  assign nw03344 = nr00001[1] ? nw03343 : nw03342;
  assign nw03345 = nr00001[2] ? nw03344 : nw03341;
  assign nw03346 = nr00001[0] ? \nr00071[25] [1] : \nr00071[24] [1];
  assign nw03347 = nr00001[0] ? \nr00071[27] [1] : \nr00071[26] [1];
  assign nw03348 = nr00001[1] ? nw03347 : nw03346;
  assign nw03349 = nr00001[0] ? \nr00071[29] [1] : \nr00071[28] [1];
  assign nw03350 = nr00001[0] ? \nr00071[31] [1] : \nr00071[30] [1];
  assign nw03351 = nr00001[1] ? nw03350 : nw03349;
  assign nw03352 = nr00001[2] ? nw03351 : nw03348;
  assign nw03353 = nr00001[3] ? nw03352 : nw03345;
  assign nw00181 = nr00001[4] ? nw03353 : nw03338;
  assign nw00328 = nw03323 ? \nr00067 [1] : nw00181;
  assign nw03354 = nr00001[0] ? \nr00071[1] [2] : \nr00071[0] [2];
  assign nw03355 = nr00001[0] ? \nr00071[3] [2] : \nr00071[2] [2];
  assign nw03356 = nr00001[1] ? nw03355 : nw03354;
  assign nw03357 = nr00001[0] ? \nr00071[5] [2] : \nr00071[4] [2];
  assign nw03358 = nr00001[0] ? \nr00071[7] [2] : \nr00071[6] [2];
  assign nw03359 = nr00001[1] ? nw03358 : nw03357;
  assign nw03360 = nr00001[2] ? nw03359 : nw03356;
  assign nw03361 = nr00001[0] ? \nr00071[9] [2] : \nr00071[8] [2];
  assign nw03362 = nr00001[0] ? \nr00071[11] [2] : \nr00071[10] [2];
  assign nw03363 = nr00001[1] ? nw03362 : nw03361;
  assign nw03364 = nr00001[0] ? \nr00071[13] [2] : \nr00071[12] [2];
  assign nw03365 = nr00001[0] ? \nr00071[15] [2] : \nr00071[14] [2];
  assign nw03366 = nr00001[1] ? nw03365 : nw03364;
  assign nw03367 = nr00001[2] ? nw03366 : nw03363;
  assign nw03368 = nr00001[3] ? nw03367 : nw03360;
  assign nw03369 = nr00001[0] ? \nr00071[17] [2] : \nr00071[16] [2];
  assign nw03370 = nr00001[0] ? \nr00071[19] [2] : \nr00071[18] [2];
  assign nw03371 = nr00001[1] ? nw03370 : nw03369;
  assign nw03372 = nr00001[0] ? \nr00071[21] [2] : \nr00071[20] [2];
  assign nw03373 = nr00001[0] ? \nr00071[23] [2] : \nr00071[22] [2];
  assign nw03374 = nr00001[1] ? nw03373 : nw03372;
  assign nw03375 = nr00001[2] ? nw03374 : nw03371;
  assign nw03376 = nr00001[0] ? \nr00071[25] [2] : \nr00071[24] [2];
  assign nw03377 = nr00001[0] ? \nr00071[27] [2] : \nr00071[26] [2];
  assign nw03378 = nr00001[1] ? nw03377 : nw03376;
  assign nw03379 = nr00001[0] ? \nr00071[29] [2] : \nr00071[28] [2];
  assign nw03380 = nr00001[0] ? \nr00071[31] [2] : \nr00071[30] [2];
  assign nw03381 = nr00001[1] ? nw03380 : nw03379;
  assign nw03382 = nr00001[2] ? nw03381 : nw03378;
  assign nw03383 = nr00001[3] ? nw03382 : nw03375;
  assign nw00192 = nr00001[4] ? nw03383 : nw03368;
  assign nw00339 = nw03323 ? \nr00067 [2] : nw00192;
  assign nw03384 = nr00001[0] ? \nr00071[1] [3] : \nr00071[0] [3];
  assign nw03385 = nr00001[0] ? \nr00071[3] [3] : \nr00071[2] [3];
  assign nw03386 = nr00001[1] ? nw03385 : nw03384;
  assign nw03387 = nr00001[0] ? \nr00071[5] [3] : \nr00071[4] [3];
  assign nw03388 = nr00001[0] ? \nr00071[7] [3] : \nr00071[6] [3];
  assign nw03389 = nr00001[1] ? nw03388 : nw03387;
  assign nw03390 = nr00001[2] ? nw03389 : nw03386;
  assign nw03391 = nr00001[0] ? \nr00071[9] [3] : \nr00071[8] [3];
  assign nw03392 = nr00001[0] ? \nr00071[11] [3] : \nr00071[10] [3];
  assign nw03393 = nr00001[1] ? nw03392 : nw03391;
  assign nw03394 = nr00001[0] ? \nr00071[13] [3] : \nr00071[12] [3];
  assign nw03395 = nr00001[0] ? \nr00071[15] [3] : \nr00071[14] [3];
  assign nw03396 = nr00001[1] ? nw03395 : nw03394;
  assign nw03397 = nr00001[2] ? nw03396 : nw03393;
  assign nw03398 = nr00001[3] ? nw03397 : nw03390;
  assign nw03399 = nr00001[0] ? \nr00071[17] [3] : \nr00071[16] [3];
  assign nw03400 = nr00001[0] ? \nr00071[19] [3] : \nr00071[18] [3];
  assign nw03401 = nr00001[1] ? nw03400 : nw03399;
  assign nw03402 = nr00001[0] ? \nr00071[21] [3] : \nr00071[20] [3];
  assign nw03403 = nr00001[0] ? \nr00071[23] [3] : \nr00071[22] [3];
  assign nw03404 = nr00001[1] ? nw03403 : nw03402;
  assign nw03405 = nr00001[2] ? nw03404 : nw03401;
  assign nw03406 = nr00001[0] ? \nr00071[25] [3] : \nr00071[24] [3];
  assign nw03407 = nr00001[0] ? \nr00071[27] [3] : \nr00071[26] [3];
  assign nw03408 = nr00001[1] ? nw03407 : nw03406;
  assign nw03409 = nr00001[0] ? \nr00071[29] [3] : \nr00071[28] [3];
  assign nw03410 = nr00001[0] ? \nr00071[31] [3] : \nr00071[30] [3];
  assign nw03411 = nr00001[1] ? nw03410 : nw03409;
  assign nw03412 = nr00001[2] ? nw03411 : nw03408;
  assign nw03413 = nr00001[3] ? nw03412 : nw03405;
  assign nw00195 = nr00001[4] ? nw03413 : nw03398;
  assign nw00342 = nw03323 ? \nr00067 [3] : nw00195;
  assign nw03414 = nr00001[0] ? \nr00071[1] [4] : \nr00071[0] [4];
  assign nw03415 = nr00001[0] ? \nr00071[3] [4] : \nr00071[2] [4];
  assign nw03416 = nr00001[1] ? nw03415 : nw03414;
  assign nw03417 = nr00001[0] ? \nr00071[5] [4] : \nr00071[4] [4];
  assign nw03418 = nr00001[0] ? \nr00071[7] [4] : \nr00071[6] [4];
  assign nw03419 = nr00001[1] ? nw03418 : nw03417;
  assign nw03420 = nr00001[2] ? nw03419 : nw03416;
  assign nw03421 = nr00001[0] ? \nr00071[9] [4] : \nr00071[8] [4];
  assign nw03422 = nr00001[0] ? \nr00071[11] [4] : \nr00071[10] [4];
  assign nw03423 = nr00001[1] ? nw03422 : nw03421;
  assign nw03424 = nr00001[0] ? \nr00071[13] [4] : \nr00071[12] [4];
  assign nw03425 = nr00001[0] ? \nr00071[15] [4] : \nr00071[14] [4];
  assign nw03426 = nr00001[1] ? nw03425 : nw03424;
  assign nw03427 = nr00001[2] ? nw03426 : nw03423;
  assign nw03428 = nr00001[3] ? nw03427 : nw03420;
  assign nw03429 = nr00001[0] ? \nr00071[17] [4] : \nr00071[16] [4];
  assign nw03430 = nr00001[0] ? \nr00071[19] [4] : \nr00071[18] [4];
  assign nw03431 = nr00001[1] ? nw03430 : nw03429;
  assign nw03432 = nr00001[0] ? \nr00071[21] [4] : \nr00071[20] [4];
  assign nw03433 = nr00001[0] ? \nr00071[23] [4] : \nr00071[22] [4];
  assign nw03434 = nr00001[1] ? nw03433 : nw03432;
  assign nw03435 = nr00001[2] ? nw03434 : nw03431;
  assign nw03436 = nr00001[0] ? \nr00071[25] [4] : \nr00071[24] [4];
  assign nw03437 = nr00001[0] ? \nr00071[27] [4] : \nr00071[26] [4];
  assign nw03438 = nr00001[1] ? nw03437 : nw03436;
  assign nw03439 = nr00001[0] ? \nr00071[29] [4] : \nr00071[28] [4];
  assign nw03440 = nr00001[0] ? \nr00071[31] [4] : \nr00071[30] [4];
  assign nw03441 = nr00001[1] ? nw03440 : nw03439;
  assign nw03442 = nr00001[2] ? nw03441 : nw03438;
  assign nw03443 = nr00001[3] ? nw03442 : nw03435;
  assign nw00196 = nr00001[4] ? nw03443 : nw03428;
  assign nw00343 = nw03323 ? \nr00067 [4] : nw00196;
  assign nw03444 = nr00001[0] ? \nr00071[1] [5] : \nr00071[0] [5];
  assign nw03445 = nr00001[0] ? \nr00071[3] [5] : \nr00071[2] [5];
  assign nw03446 = nr00001[1] ? nw03445 : nw03444;
  assign nw03447 = nr00001[0] ? \nr00071[5] [5] : \nr00071[4] [5];
  assign nw03448 = nr00001[0] ? \nr00071[7] [5] : \nr00071[6] [5];
  assign nw03449 = nr00001[1] ? nw03448 : nw03447;
  assign nw03450 = nr00001[2] ? nw03449 : nw03446;
  assign nw03451 = nr00001[0] ? \nr00071[9] [5] : \nr00071[8] [5];
  assign nw03452 = nr00001[0] ? \nr00071[11] [5] : \nr00071[10] [5];
  assign nw03453 = nr00001[1] ? nw03452 : nw03451;
  assign nw03454 = nr00001[0] ? \nr00071[13] [5] : \nr00071[12] [5];
  assign nw03455 = nr00001[0] ? \nr00071[15] [5] : \nr00071[14] [5];
  assign nw03456 = nr00001[1] ? nw03455 : nw03454;
  assign nw03457 = nr00001[2] ? nw03456 : nw03453;
  assign nw03458 = nr00001[3] ? nw03457 : nw03450;
  assign nw03459 = nr00001[0] ? \nr00071[17] [5] : \nr00071[16] [5];
  assign nw03460 = nr00001[0] ? \nr00071[19] [5] : \nr00071[18] [5];
  assign nw03461 = nr00001[1] ? nw03460 : nw03459;
  assign nw03462 = nr00001[0] ? \nr00071[21] [5] : \nr00071[20] [5];
  assign nw03463 = nr00001[0] ? \nr00071[23] [5] : \nr00071[22] [5];
  assign nw03464 = nr00001[1] ? nw03463 : nw03462;
  assign nw03465 = nr00001[2] ? nw03464 : nw03461;
  assign nw03466 = nr00001[0] ? \nr00071[25] [5] : \nr00071[24] [5];
  assign nw03467 = nr00001[0] ? \nr00071[27] [5] : \nr00071[26] [5];
  assign nw03468 = nr00001[1] ? nw03467 : nw03466;
  assign nw03469 = nr00001[0] ? \nr00071[29] [5] : \nr00071[28] [5];
  assign nw03470 = nr00001[0] ? \nr00071[31] [5] : \nr00071[30] [5];
  assign nw03471 = nr00001[1] ? nw03470 : nw03469;
  assign nw03472 = nr00001[2] ? nw03471 : nw03468;
  assign nw03473 = nr00001[3] ? nw03472 : nw03465;
  assign nw00197 = nr00001[4] ? nw03473 : nw03458;
  assign nw00344 = nw03323 ? \nr00067 [5] : nw00197;
  assign nw03474 = nr00001[0] ? \nr00071[1] [6] : \nr00071[0] [6];
  assign nw03475 = nr00001[0] ? \nr00071[3] [6] : \nr00071[2] [6];
  assign nw03476 = nr00001[1] ? nw03475 : nw03474;
  assign nw03477 = nr00001[0] ? \nr00071[5] [6] : \nr00071[4] [6];
  assign nw03478 = nr00001[0] ? \nr00071[7] [6] : \nr00071[6] [6];
  assign nw03479 = nr00001[1] ? nw03478 : nw03477;
  assign nw03480 = nr00001[2] ? nw03479 : nw03476;
  assign nw03481 = nr00001[0] ? \nr00071[9] [6] : \nr00071[8] [6];
  assign nw03482 = nr00001[0] ? \nr00071[11] [6] : \nr00071[10] [6];
  assign nw03483 = nr00001[1] ? nw03482 : nw03481;
  assign nw03484 = nr00001[0] ? \nr00071[13] [6] : \nr00071[12] [6];
  assign nw03485 = nr00001[0] ? \nr00071[15] [6] : \nr00071[14] [6];
  assign nw03486 = nr00001[1] ? nw03485 : nw03484;
  assign nw03487 = nr00001[2] ? nw03486 : nw03483;
  assign nw03488 = nr00001[3] ? nw03487 : nw03480;
  assign nw03489 = nr00001[0] ? \nr00071[17] [6] : \nr00071[16] [6];
  assign nw03490 = nr00001[0] ? \nr00071[19] [6] : \nr00071[18] [6];
  assign nw03491 = nr00001[1] ? nw03490 : nw03489;
  assign nw03492 = nr00001[0] ? \nr00071[21] [6] : \nr00071[20] [6];
  assign nw03493 = nr00001[0] ? \nr00071[23] [6] : \nr00071[22] [6];
  assign nw03494 = nr00001[1] ? nw03493 : nw03492;
  assign nw03495 = nr00001[2] ? nw03494 : nw03491;
  assign nw03496 = nr00001[0] ? \nr00071[25] [6] : \nr00071[24] [6];
  assign nw03497 = nr00001[0] ? \nr00071[27] [6] : \nr00071[26] [6];
  assign nw03498 = nr00001[1] ? nw03497 : nw03496;
  assign nw03499 = nr00001[0] ? \nr00071[29] [6] : \nr00071[28] [6];
  assign nw03500 = nr00001[0] ? \nr00071[31] [6] : \nr00071[30] [6];
  assign nw03501 = nr00001[1] ? nw03500 : nw03499;
  assign nw03502 = nr00001[2] ? nw03501 : nw03498;
  assign nw03503 = nr00001[3] ? nw03502 : nw03495;
  assign nw00198 = nr00001[4] ? nw03503 : nw03488;
  assign nw00345 = nw03323 ? \nr00067 [6] : nw00198;
  assign nw03504 = nr00001[0] ? \nr00071[1] [7] : \nr00071[0] [7];
  assign nw03505 = nr00001[0] ? \nr00071[3] [7] : \nr00071[2] [7];
  assign nw03506 = nr00001[1] ? nw03505 : nw03504;
  assign nw03507 = nr00001[0] ? \nr00071[5] [7] : \nr00071[4] [7];
  assign nw03508 = nr00001[0] ? \nr00071[7] [7] : \nr00071[6] [7];
  assign nw03509 = nr00001[1] ? nw03508 : nw03507;
  assign nw03510 = nr00001[2] ? nw03509 : nw03506;
  assign nw03511 = nr00001[0] ? \nr00071[9] [7] : \nr00071[8] [7];
  assign nw03512 = nr00001[0] ? \nr00071[11] [7] : \nr00071[10] [7];
  assign nw03513 = nr00001[1] ? nw03512 : nw03511;
  assign nw03514 = nr00001[0] ? \nr00071[13] [7] : \nr00071[12] [7];
  assign nw03515 = nr00001[0] ? \nr00071[15] [7] : \nr00071[14] [7];
  assign nw03516 = nr00001[1] ? nw03515 : nw03514;
  assign nw03517 = nr00001[2] ? nw03516 : nw03513;
  assign nw03518 = nr00001[3] ? nw03517 : nw03510;
  assign nw03519 = nr00001[0] ? \nr00071[17] [7] : \nr00071[16] [7];
  assign nw03520 = nr00001[0] ? \nr00071[19] [7] : \nr00071[18] [7];
  assign nw03521 = nr00001[1] ? nw03520 : nw03519;
  assign nw03522 = nr00001[0] ? \nr00071[21] [7] : \nr00071[20] [7];
  assign nw03523 = nr00001[0] ? \nr00071[23] [7] : \nr00071[22] [7];
  assign nw03524 = nr00001[1] ? nw03523 : nw03522;
  assign nw03525 = nr00001[2] ? nw03524 : nw03521;
  assign nw03526 = nr00001[0] ? \nr00071[25] [7] : \nr00071[24] [7];
  assign nw03527 = nr00001[0] ? \nr00071[27] [7] : \nr00071[26] [7];
  assign nw03528 = nr00001[1] ? nw03527 : nw03526;
  assign nw03529 = nr00001[0] ? \nr00071[29] [7] : \nr00071[28] [7];
  assign nw03530 = nr00001[0] ? \nr00071[31] [7] : \nr00071[30] [7];
  assign nw03531 = nr00001[1] ? nw03530 : nw03529;
  assign nw03532 = nr00001[2] ? nw03531 : nw03528;
  assign nw03533 = nr00001[3] ? nw03532 : nw03525;
  assign nw00199 = nr00001[4] ? nw03533 : nw03518;
  assign nw00346 = nw03323 ? \nr00067 [7] : nw00199;
  assign nw03534 = nr00001[0] ? \nr00071[1] [8] : \nr00071[0] [8];
  assign nw03535 = nr00001[0] ? \nr00071[3] [8] : \nr00071[2] [8];
  assign nw03536 = nr00001[1] ? nw03535 : nw03534;
  assign nw03537 = nr00001[0] ? \nr00071[5] [8] : \nr00071[4] [8];
  assign nw03538 = nr00001[0] ? \nr00071[7] [8] : \nr00071[6] [8];
  assign nw03539 = nr00001[1] ? nw03538 : nw03537;
  assign nw03540 = nr00001[2] ? nw03539 : nw03536;
  assign nw03541 = nr00001[0] ? \nr00071[9] [8] : \nr00071[8] [8];
  assign nw03542 = nr00001[0] ? \nr00071[11] [8] : \nr00071[10] [8];
  assign nw03543 = nr00001[1] ? nw03542 : nw03541;
  assign nw03544 = nr00001[0] ? \nr00071[13] [8] : \nr00071[12] [8];
  assign nw03545 = nr00001[0] ? \nr00071[15] [8] : \nr00071[14] [8];
  assign nw03546 = nr00001[1] ? nw03545 : nw03544;
  assign nw03547 = nr00001[2] ? nw03546 : nw03543;
  assign nw03548 = nr00001[3] ? nw03547 : nw03540;
  assign nw03549 = nr00001[0] ? \nr00071[17] [8] : \nr00071[16] [8];
  assign nw03550 = nr00001[0] ? \nr00071[19] [8] : \nr00071[18] [8];
  assign nw03551 = nr00001[1] ? nw03550 : nw03549;
  assign nw03552 = nr00001[0] ? \nr00071[21] [8] : \nr00071[20] [8];
  assign nw03553 = nr00001[0] ? \nr00071[23] [8] : \nr00071[22] [8];
  assign nw03554 = nr00001[1] ? nw03553 : nw03552;
  assign nw03555 = nr00001[2] ? nw03554 : nw03551;
  assign nw03556 = nr00001[0] ? \nr00071[25] [8] : \nr00071[24] [8];
  assign nw03557 = nr00001[0] ? \nr00071[27] [8] : \nr00071[26] [8];
  assign nw03558 = nr00001[1] ? nw03557 : nw03556;
  assign nw03559 = nr00001[0] ? \nr00071[29] [8] : \nr00071[28] [8];
  assign nw03560 = nr00001[0] ? \nr00071[31] [8] : \nr00071[30] [8];
  assign nw03561 = nr00001[1] ? nw03560 : nw03559;
  assign nw03562 = nr00001[2] ? nw03561 : nw03558;
  assign nw03563 = nr00001[3] ? nw03562 : nw03555;
  assign nw00200 = nr00001[4] ? nw03563 : nw03548;
  assign nw00347 = nw03323 ? \nr00067 [8] : nw00200;
  assign nw03564 = nr00001[0] ? \nr00071[1] [9] : \nr00071[0] [9];
  assign nw03565 = nr00001[0] ? \nr00071[3] [9] : \nr00071[2] [9];
  assign nw03566 = nr00001[1] ? nw03565 : nw03564;
  assign nw03567 = nr00001[0] ? \nr00071[5] [9] : \nr00071[4] [9];
  assign nw03568 = nr00001[0] ? \nr00071[7] [9] : \nr00071[6] [9];
  assign nw03569 = nr00001[1] ? nw03568 : nw03567;
  assign nw03570 = nr00001[2] ? nw03569 : nw03566;
  assign nw03571 = nr00001[0] ? \nr00071[9] [9] : \nr00071[8] [9];
  assign nw03572 = nr00001[0] ? \nr00071[11] [9] : \nr00071[10] [9];
  assign nw03573 = nr00001[1] ? nw03572 : nw03571;
  assign nw03574 = nr00001[0] ? \nr00071[13] [9] : \nr00071[12] [9];
  assign nw03575 = nr00001[0] ? \nr00071[15] [9] : \nr00071[14] [9];
  assign nw03576 = nr00001[1] ? nw03575 : nw03574;
  assign nw03577 = nr00001[2] ? nw03576 : nw03573;
  assign nw03578 = nr00001[3] ? nw03577 : nw03570;
  assign nw03579 = nr00001[0] ? \nr00071[17] [9] : \nr00071[16] [9];
  assign nw03580 = nr00001[0] ? \nr00071[19] [9] : \nr00071[18] [9];
  assign nw03581 = nr00001[1] ? nw03580 : nw03579;
  assign nw03582 = nr00001[0] ? \nr00071[21] [9] : \nr00071[20] [9];
  assign nw03583 = nr00001[0] ? \nr00071[23] [9] : \nr00071[22] [9];
  assign nw03584 = nr00001[1] ? nw03583 : nw03582;
  assign nw03585 = nr00001[2] ? nw03584 : nw03581;
  assign nw03586 = nr00001[0] ? \nr00071[25] [9] : \nr00071[24] [9];
  assign nw03587 = nr00001[0] ? \nr00071[27] [9] : \nr00071[26] [9];
  assign nw03588 = nr00001[1] ? nw03587 : nw03586;
  assign nw03589 = nr00001[0] ? \nr00071[29] [9] : \nr00071[28] [9];
  assign nw03590 = nr00001[0] ? \nr00071[31] [9] : \nr00071[30] [9];
  assign nw03591 = nr00001[1] ? nw03590 : nw03589;
  assign nw03592 = nr00001[2] ? nw03591 : nw03588;
  assign nw03593 = nr00001[3] ? nw03592 : nw03585;
  assign nw00201 = nr00001[4] ? nw03593 : nw03578;
  assign nw00348 = nw03323 ? \nr00067 [9] : nw00201;
  assign nw03594 = nr00001[0] ? \nr00071[1] [10] : \nr00071[0] [10];
  assign nw03595 = nr00001[0] ? \nr00071[3] [10] : \nr00071[2] [10];
  assign nw03596 = nr00001[1] ? nw03595 : nw03594;
  assign nw03597 = nr00001[0] ? \nr00071[5] [10] : \nr00071[4] [10];
  assign nw03598 = nr00001[0] ? \nr00071[7] [10] : \nr00071[6] [10];
  assign nw03599 = nr00001[1] ? nw03598 : nw03597;
  assign nw03600 = nr00001[2] ? nw03599 : nw03596;
  assign nw03601 = nr00001[0] ? \nr00071[9] [10] : \nr00071[8] [10];
  assign nw03602 = nr00001[0] ? \nr00071[11] [10] : \nr00071[10] [10];
  assign nw03603 = nr00001[1] ? nw03602 : nw03601;
  assign nw03604 = nr00001[0] ? \nr00071[13] [10] : \nr00071[12] [10];
  assign nw03605 = nr00001[0] ? \nr00071[15] [10] : \nr00071[14] [10];
  assign nw03606 = nr00001[1] ? nw03605 : nw03604;
  assign nw03607 = nr00001[2] ? nw03606 : nw03603;
  assign nw03608 = nr00001[3] ? nw03607 : nw03600;
  assign nw03609 = nr00001[0] ? \nr00071[17] [10] : \nr00071[16] [10];
  assign nw03610 = nr00001[0] ? \nr00071[19] [10] : \nr00071[18] [10];
  assign nw03611 = nr00001[1] ? nw03610 : nw03609;
  assign nw03612 = nr00001[0] ? \nr00071[21] [10] : \nr00071[20] [10];
  assign nw03613 = nr00001[0] ? \nr00071[23] [10] : \nr00071[22] [10];
  assign nw03614 = nr00001[1] ? nw03613 : nw03612;
  assign nw03615 = nr00001[2] ? nw03614 : nw03611;
  assign nw03616 = nr00001[0] ? \nr00071[25] [10] : \nr00071[24] [10];
  assign nw03617 = nr00001[0] ? \nr00071[27] [10] : \nr00071[26] [10];
  assign nw03618 = nr00001[1] ? nw03617 : nw03616;
  assign nw03619 = nr00001[0] ? \nr00071[29] [10] : \nr00071[28] [10];
  assign nw03620 = nr00001[0] ? \nr00071[31] [10] : \nr00071[30] [10];
  assign nw03621 = nr00001[1] ? nw03620 : nw03619;
  assign nw03622 = nr00001[2] ? nw03621 : nw03618;
  assign nw03623 = nr00001[3] ? nw03622 : nw03615;
  assign nw00171 = nr00001[4] ? nw03623 : nw03608;
  assign nw00318 = nw03323 ? \nr00067 [10] : nw00171;
  assign nw03624 = nr00001[0] ? \nr00071[1] [11] : \nr00071[0] [11];
  assign nw03625 = nr00001[0] ? \nr00071[3] [11] : \nr00071[2] [11];
  assign nw03626 = nr00001[1] ? nw03625 : nw03624;
  assign nw03627 = nr00001[0] ? \nr00071[5] [11] : \nr00071[4] [11];
  assign nw03628 = nr00001[0] ? \nr00071[7] [11] : \nr00071[6] [11];
  assign nw03629 = nr00001[1] ? nw03628 : nw03627;
  assign nw03630 = nr00001[2] ? nw03629 : nw03626;
  assign nw03631 = nr00001[0] ? \nr00071[9] [11] : \nr00071[8] [11];
  assign nw03632 = nr00001[0] ? \nr00071[11] [11] : \nr00071[10] [11];
  assign nw03633 = nr00001[1] ? nw03632 : nw03631;
  assign nw03634 = nr00001[0] ? \nr00071[13] [11] : \nr00071[12] [11];
  assign nw03635 = nr00001[0] ? \nr00071[15] [11] : \nr00071[14] [11];
  assign nw03636 = nr00001[1] ? nw03635 : nw03634;
  assign nw03637 = nr00001[2] ? nw03636 : nw03633;
  assign nw03638 = nr00001[3] ? nw03637 : nw03630;
  assign nw03639 = nr00001[0] ? \nr00071[17] [11] : \nr00071[16] [11];
  assign nw03640 = nr00001[0] ? \nr00071[19] [11] : \nr00071[18] [11];
  assign nw03641 = nr00001[1] ? nw03640 : nw03639;
  assign nw03642 = nr00001[0] ? \nr00071[21] [11] : \nr00071[20] [11];
  assign nw03643 = nr00001[0] ? \nr00071[23] [11] : \nr00071[22] [11];
  assign nw03644 = nr00001[1] ? nw03643 : nw03642;
  assign nw03645 = nr00001[2] ? nw03644 : nw03641;
  assign nw03646 = nr00001[0] ? \nr00071[25] [11] : \nr00071[24] [11];
  assign nw03647 = nr00001[0] ? \nr00071[27] [11] : \nr00071[26] [11];
  assign nw03648 = nr00001[1] ? nw03647 : nw03646;
  assign nw03649 = nr00001[0] ? \nr00071[29] [11] : \nr00071[28] [11];
  assign nw03650 = nr00001[0] ? \nr00071[31] [11] : \nr00071[30] [11];
  assign nw03651 = nr00001[1] ? nw03650 : nw03649;
  assign nw03652 = nr00001[2] ? nw03651 : nw03648;
  assign nw03653 = nr00001[3] ? nw03652 : nw03645;
  assign nw00172 = nr00001[4] ? nw03653 : nw03638;
  assign nw00319 = nw03323 ? \nr00067 [11] : nw00172;
  assign nw03654 = nr00001[0] ? \nr00071[1] [12] : \nr00071[0] [12];
  assign nw03655 = nr00001[0] ? \nr00071[3] [12] : \nr00071[2] [12];
  assign nw03656 = nr00001[1] ? nw03655 : nw03654;
  assign nw03657 = nr00001[0] ? \nr00071[5] [12] : \nr00071[4] [12];
  assign nw03658 = nr00001[0] ? \nr00071[7] [12] : \nr00071[6] [12];
  assign nw03659 = nr00001[1] ? nw03658 : nw03657;
  assign nw03660 = nr00001[2] ? nw03659 : nw03656;
  assign nw03661 = nr00001[0] ? \nr00071[9] [12] : \nr00071[8] [12];
  assign nw03662 = nr00001[0] ? \nr00071[11] [12] : \nr00071[10] [12];
  assign nw03663 = nr00001[1] ? nw03662 : nw03661;
  assign nw03664 = nr00001[0] ? \nr00071[13] [12] : \nr00071[12] [12];
  assign nw03665 = nr00001[0] ? \nr00071[15] [12] : \nr00071[14] [12];
  assign nw03666 = nr00001[1] ? nw03665 : nw03664;
  assign nw03667 = nr00001[2] ? nw03666 : nw03663;
  assign nw03668 = nr00001[3] ? nw03667 : nw03660;
  assign nw03669 = nr00001[0] ? \nr00071[17] [12] : \nr00071[16] [12];
  assign nw03670 = nr00001[0] ? \nr00071[19] [12] : \nr00071[18] [12];
  assign nw03671 = nr00001[1] ? nw03670 : nw03669;
  assign nw03672 = nr00001[0] ? \nr00071[21] [12] : \nr00071[20] [12];
  assign nw03673 = nr00001[0] ? \nr00071[23] [12] : \nr00071[22] [12];
  assign nw03674 = nr00001[1] ? nw03673 : nw03672;
  assign nw03675 = nr00001[2] ? nw03674 : nw03671;
  assign nw03676 = nr00001[0] ? \nr00071[25] [12] : \nr00071[24] [12];
  assign nw03677 = nr00001[0] ? \nr00071[27] [12] : \nr00071[26] [12];
  assign nw03678 = nr00001[1] ? nw03677 : nw03676;
  assign nw03679 = nr00001[0] ? \nr00071[29] [12] : \nr00071[28] [12];
  assign nw03680 = nr00001[0] ? \nr00071[31] [12] : \nr00071[30] [12];
  assign nw03681 = nr00001[1] ? nw03680 : nw03679;
  assign nw03682 = nr00001[2] ? nw03681 : nw03678;
  assign nw03683 = nr00001[3] ? nw03682 : nw03675;
  assign nw00173 = nr00001[4] ? nw03683 : nw03668;
  assign nw00320 = nw03323 ? \nr00067 [12] : nw00173;
  assign nw03684 = nr00001[0] ? \nr00071[1] [13] : \nr00071[0] [13];
  assign nw03685 = nr00001[0] ? \nr00071[3] [13] : \nr00071[2] [13];
  assign nw03686 = nr00001[1] ? nw03685 : nw03684;
  assign nw03687 = nr00001[0] ? \nr00071[5] [13] : \nr00071[4] [13];
  assign nw03688 = nr00001[0] ? \nr00071[7] [13] : \nr00071[6] [13];
  assign nw03689 = nr00001[1] ? nw03688 : nw03687;
  assign nw03690 = nr00001[2] ? nw03689 : nw03686;
  assign nw03691 = nr00001[0] ? \nr00071[9] [13] : \nr00071[8] [13];
  assign nw03692 = nr00001[0] ? \nr00071[11] [13] : \nr00071[10] [13];
  assign nw03693 = nr00001[1] ? nw03692 : nw03691;
  assign nw03694 = nr00001[0] ? \nr00071[13] [13] : \nr00071[12] [13];
  assign nw03695 = nr00001[0] ? \nr00071[15] [13] : \nr00071[14] [13];
  assign nw03696 = nr00001[1] ? nw03695 : nw03694;
  assign nw03697 = nr00001[2] ? nw03696 : nw03693;
  assign nw03698 = nr00001[3] ? nw03697 : nw03690;
  assign nw03699 = nr00001[0] ? \nr00071[17] [13] : \nr00071[16] [13];
  assign nw03700 = nr00001[0] ? \nr00071[19] [13] : \nr00071[18] [13];
  assign nw03701 = nr00001[1] ? nw03700 : nw03699;
  assign nw03702 = nr00001[0] ? \nr00071[21] [13] : \nr00071[20] [13];
  assign nw03703 = nr00001[0] ? \nr00071[23] [13] : \nr00071[22] [13];
  assign nw03704 = nr00001[1] ? nw03703 : nw03702;
  assign nw03705 = nr00001[2] ? nw03704 : nw03701;
  assign nw03706 = nr00001[0] ? \nr00071[25] [13] : \nr00071[24] [13];
  assign nw03707 = nr00001[0] ? \nr00071[27] [13] : \nr00071[26] [13];
  assign nw03708 = nr00001[1] ? nw03707 : nw03706;
  assign nw03709 = nr00001[0] ? \nr00071[29] [13] : \nr00071[28] [13];
  assign nw03710 = nr00001[0] ? \nr00071[31] [13] : \nr00071[30] [13];
  assign nw03711 = nr00001[1] ? nw03710 : nw03709;
  assign nw03712 = nr00001[2] ? nw03711 : nw03708;
  assign nw03713 = nr00001[3] ? nw03712 : nw03705;
  assign nw00174 = nr00001[4] ? nw03713 : nw03698;
  assign nw00321 = nw03323 ? \nr00067 [13] : nw00174;
  assign nw03714 = nr00001[0] ? \nr00071[1] [14] : \nr00071[0] [14];
  assign nw03715 = nr00001[0] ? \nr00071[3] [14] : \nr00071[2] [14];
  assign nw03716 = nr00001[1] ? nw03715 : nw03714;
  assign nw03717 = nr00001[0] ? \nr00071[5] [14] : \nr00071[4] [14];
  assign nw03718 = nr00001[0] ? \nr00071[7] [14] : \nr00071[6] [14];
  assign nw03719 = nr00001[1] ? nw03718 : nw03717;
  assign nw03720 = nr00001[2] ? nw03719 : nw03716;
  assign nw03721 = nr00001[0] ? \nr00071[9] [14] : \nr00071[8] [14];
  assign nw03722 = nr00001[0] ? \nr00071[11] [14] : \nr00071[10] [14];
  assign nw03723 = nr00001[1] ? nw03722 : nw03721;
  assign nw03724 = nr00001[0] ? \nr00071[13] [14] : \nr00071[12] [14];
  assign nw03725 = nr00001[0] ? \nr00071[15] [14] : \nr00071[14] [14];
  assign nw03726 = nr00001[1] ? nw03725 : nw03724;
  assign nw03727 = nr00001[2] ? nw03726 : nw03723;
  assign nw03728 = nr00001[3] ? nw03727 : nw03720;
  assign nw03729 = nr00001[0] ? \nr00071[17] [14] : \nr00071[16] [14];
  assign nw03730 = nr00001[0] ? \nr00071[19] [14] : \nr00071[18] [14];
  assign nw03731 = nr00001[1] ? nw03730 : nw03729;
  assign nw03732 = nr00001[0] ? \nr00071[21] [14] : \nr00071[20] [14];
  assign nw03733 = nr00001[0] ? \nr00071[23] [14] : \nr00071[22] [14];
  assign nw03734 = nr00001[1] ? nw03733 : nw03732;
  assign nw03735 = nr00001[2] ? nw03734 : nw03731;
  assign nw03736 = nr00001[0] ? \nr00071[25] [14] : \nr00071[24] [14];
  assign nw03737 = nr00001[0] ? \nr00071[27] [14] : \nr00071[26] [14];
  assign nw03738 = nr00001[1] ? nw03737 : nw03736;
  assign nw03739 = nr00001[0] ? \nr00071[29] [14] : \nr00071[28] [14];
  assign nw03740 = nr00001[0] ? \nr00071[31] [14] : \nr00071[30] [14];
  assign nw03741 = nr00001[1] ? nw03740 : nw03739;
  assign nw03742 = nr00001[2] ? nw03741 : nw03738;
  assign nw03743 = nr00001[3] ? nw03742 : nw03735;
  assign nw00175 = nr00001[4] ? nw03743 : nw03728;
  assign nw00322 = nw03323 ? \nr00067 [14] : nw00175;
  assign nw03744 = nr00001[0] ? \nr00071[1] [15] : \nr00071[0] [15];
  assign nw03745 = nr00001[0] ? \nr00071[3] [15] : \nr00071[2] [15];
  assign nw03746 = nr00001[1] ? nw03745 : nw03744;
  assign nw03747 = nr00001[0] ? \nr00071[5] [15] : \nr00071[4] [15];
  assign nw03748 = nr00001[0] ? \nr00071[7] [15] : \nr00071[6] [15];
  assign nw03749 = nr00001[1] ? nw03748 : nw03747;
  assign nw03750 = nr00001[2] ? nw03749 : nw03746;
  assign nw03751 = nr00001[0] ? \nr00071[9] [15] : \nr00071[8] [15];
  assign nw03752 = nr00001[0] ? \nr00071[11] [15] : \nr00071[10] [15];
  assign nw03753 = nr00001[1] ? nw03752 : nw03751;
  assign nw03754 = nr00001[0] ? \nr00071[13] [15] : \nr00071[12] [15];
  assign nw03755 = nr00001[0] ? \nr00071[15] [15] : \nr00071[14] [15];
  assign nw03756 = nr00001[1] ? nw03755 : nw03754;
  assign nw03757 = nr00001[2] ? nw03756 : nw03753;
  assign nw03758 = nr00001[3] ? nw03757 : nw03750;
  assign nw03759 = nr00001[0] ? \nr00071[17] [15] : \nr00071[16] [15];
  assign nw03760 = nr00001[0] ? \nr00071[19] [15] : \nr00071[18] [15];
  assign nw03761 = nr00001[1] ? nw03760 : nw03759;
  assign nw03762 = nr00001[0] ? \nr00071[21] [15] : \nr00071[20] [15];
  assign nw03763 = nr00001[0] ? \nr00071[23] [15] : \nr00071[22] [15];
  assign nw03764 = nr00001[1] ? nw03763 : nw03762;
  assign nw03765 = nr00001[2] ? nw03764 : nw03761;
  assign nw03766 = nr00001[0] ? \nr00071[25] [15] : \nr00071[24] [15];
  assign nw03767 = nr00001[0] ? \nr00071[27] [15] : \nr00071[26] [15];
  assign nw03768 = nr00001[1] ? nw03767 : nw03766;
  assign nw03769 = nr00001[0] ? \nr00071[29] [15] : \nr00071[28] [15];
  assign nw03770 = nr00001[0] ? \nr00071[31] [15] : \nr00071[30] [15];
  assign nw03771 = nr00001[1] ? nw03770 : nw03769;
  assign nw03772 = nr00001[2] ? nw03771 : nw03768;
  assign nw03773 = nr00001[3] ? nw03772 : nw03765;
  assign nw00176 = nr00001[4] ? nw03773 : nw03758;
  assign nw00323 = nw03323 ? \nr00067 [15] : nw00176;
  assign nw03774 = nr00001[0] ? \nr00071[1] [16] : \nr00071[0] [16];
  assign nw03775 = nr00001[0] ? \nr00071[3] [16] : \nr00071[2] [16];
  assign nw03776 = nr00001[1] ? nw03775 : nw03774;
  assign nw03777 = nr00001[0] ? \nr00071[5] [16] : \nr00071[4] [16];
  assign nw03778 = nr00001[0] ? \nr00071[7] [16] : \nr00071[6] [16];
  assign nw03779 = nr00001[1] ? nw03778 : nw03777;
  assign nw03780 = nr00001[2] ? nw03779 : nw03776;
  assign nw03781 = nr00001[0] ? \nr00071[9] [16] : \nr00071[8] [16];
  assign nw03782 = nr00001[0] ? \nr00071[11] [16] : \nr00071[10] [16];
  assign nw03783 = nr00001[1] ? nw03782 : nw03781;
  assign nw03784 = nr00001[0] ? \nr00071[13] [16] : \nr00071[12] [16];
  assign nw03785 = nr00001[0] ? \nr00071[15] [16] : \nr00071[14] [16];
  assign nw03786 = nr00001[1] ? nw03785 : nw03784;
  assign nw03787 = nr00001[2] ? nw03786 : nw03783;
  assign nw03788 = nr00001[3] ? nw03787 : nw03780;
  assign nw03789 = nr00001[0] ? \nr00071[17] [16] : \nr00071[16] [16];
  assign nw03790 = nr00001[0] ? \nr00071[19] [16] : \nr00071[18] [16];
  assign nw03791 = nr00001[1] ? nw03790 : nw03789;
  assign nw03792 = nr00001[0] ? \nr00071[21] [16] : \nr00071[20] [16];
  assign nw03793 = nr00001[0] ? \nr00071[23] [16] : \nr00071[22] [16];
  assign nw03794 = nr00001[1] ? nw03793 : nw03792;
  assign nw03795 = nr00001[2] ? nw03794 : nw03791;
  assign nw03796 = nr00001[0] ? \nr00071[25] [16] : \nr00071[24] [16];
  assign nw03797 = nr00001[0] ? \nr00071[27] [16] : \nr00071[26] [16];
  assign nw03798 = nr00001[1] ? nw03797 : nw03796;
  assign nw03799 = nr00001[0] ? \nr00071[29] [16] : \nr00071[28] [16];
  assign nw03800 = nr00001[0] ? \nr00071[31] [16] : \nr00071[30] [16];
  assign nw03801 = nr00001[1] ? nw03800 : nw03799;
  assign nw03802 = nr00001[2] ? nw03801 : nw03798;
  assign nw03803 = nr00001[3] ? nw03802 : nw03795;
  assign nw00177 = nr00001[4] ? nw03803 : nw03788;
  assign nw00324 = nw03323 ? \nr00067 [16] : nw00177;
  assign nw03804 = nr00001[0] ? \nr00071[1] [17] : \nr00071[0] [17];
  assign nw03805 = nr00001[0] ? \nr00071[3] [17] : \nr00071[2] [17];
  assign nw03806 = nr00001[1] ? nw03805 : nw03804;
  assign nw03807 = nr00001[0] ? \nr00071[5] [17] : \nr00071[4] [17];
  assign nw03808 = nr00001[0] ? \nr00071[7] [17] : \nr00071[6] [17];
  assign nw03809 = nr00001[1] ? nw03808 : nw03807;
  assign nw03810 = nr00001[2] ? nw03809 : nw03806;
  assign nw03811 = nr00001[0] ? \nr00071[9] [17] : \nr00071[8] [17];
  assign nw03812 = nr00001[0] ? \nr00071[11] [17] : \nr00071[10] [17];
  assign nw03813 = nr00001[1] ? nw03812 : nw03811;
  assign nw03814 = nr00001[0] ? \nr00071[13] [17] : \nr00071[12] [17];
  assign nw03815 = nr00001[0] ? \nr00071[15] [17] : \nr00071[14] [17];
  assign nw03816 = nr00001[1] ? nw03815 : nw03814;
  assign nw03817 = nr00001[2] ? nw03816 : nw03813;
  assign nw03818 = nr00001[3] ? nw03817 : nw03810;
  assign nw03819 = nr00001[0] ? \nr00071[17] [17] : \nr00071[16] [17];
  assign nw03820 = nr00001[0] ? \nr00071[19] [17] : \nr00071[18] [17];
  assign nw03821 = nr00001[1] ? nw03820 : nw03819;
  assign nw03822 = nr00001[0] ? \nr00071[21] [17] : \nr00071[20] [17];
  assign nw03823 = nr00001[0] ? \nr00071[23] [17] : \nr00071[22] [17];
  assign nw03824 = nr00001[1] ? nw03823 : nw03822;
  assign nw03825 = nr00001[2] ? nw03824 : nw03821;
  assign nw03826 = nr00001[0] ? \nr00071[25] [17] : \nr00071[24] [17];
  assign nw03827 = nr00001[0] ? \nr00071[27] [17] : \nr00071[26] [17];
  assign nw03828 = nr00001[1] ? nw03827 : nw03826;
  assign nw03829 = nr00001[0] ? \nr00071[29] [17] : \nr00071[28] [17];
  assign nw03830 = nr00001[0] ? \nr00071[31] [17] : \nr00071[30] [17];
  assign nw03831 = nr00001[1] ? nw03830 : nw03829;
  assign nw03832 = nr00001[2] ? nw03831 : nw03828;
  assign nw03833 = nr00001[3] ? nw03832 : nw03825;
  assign nw00178 = nr00001[4] ? nw03833 : nw03818;
  assign nw00325 = nw03323 ? \nr00067 [17] : nw00178;
  assign nw03834 = nr00001[0] ? \nr00071[1] [18] : \nr00071[0] [18];
  assign nw03835 = nr00001[0] ? \nr00071[3] [18] : \nr00071[2] [18];
  assign nw03836 = nr00001[1] ? nw03835 : nw03834;
  assign nw03837 = nr00001[0] ? \nr00071[5] [18] : \nr00071[4] [18];
  assign nw03838 = nr00001[0] ? \nr00071[7] [18] : \nr00071[6] [18];
  assign nw03839 = nr00001[1] ? nw03838 : nw03837;
  assign nw03840 = nr00001[2] ? nw03839 : nw03836;
  assign nw03841 = nr00001[0] ? \nr00071[9] [18] : \nr00071[8] [18];
  assign nw03842 = nr00001[0] ? \nr00071[11] [18] : \nr00071[10] [18];
  assign nw03843 = nr00001[1] ? nw03842 : nw03841;
  assign nw03844 = nr00001[0] ? \nr00071[13] [18] : \nr00071[12] [18];
  assign nw03845 = nr00001[0] ? \nr00071[15] [18] : \nr00071[14] [18];
  assign nw03846 = nr00001[1] ? nw03845 : nw03844;
  assign nw03847 = nr00001[2] ? nw03846 : nw03843;
  assign nw03848 = nr00001[3] ? nw03847 : nw03840;
  assign nw03849 = nr00001[0] ? \nr00071[17] [18] : \nr00071[16] [18];
  assign nw03850 = nr00001[0] ? \nr00071[19] [18] : \nr00071[18] [18];
  assign nw03851 = nr00001[1] ? nw03850 : nw03849;
  assign nw03852 = nr00001[0] ? \nr00071[21] [18] : \nr00071[20] [18];
  assign nw03853 = nr00001[0] ? \nr00071[23] [18] : \nr00071[22] [18];
  assign nw03854 = nr00001[1] ? nw03853 : nw03852;
  assign nw03855 = nr00001[2] ? nw03854 : nw03851;
  assign nw03856 = nr00001[0] ? \nr00071[25] [18] : \nr00071[24] [18];
  assign nw03857 = nr00001[0] ? \nr00071[27] [18] : \nr00071[26] [18];
  assign nw03858 = nr00001[1] ? nw03857 : nw03856;
  assign nw03859 = nr00001[0] ? \nr00071[29] [18] : \nr00071[28] [18];
  assign nw03860 = nr00001[0] ? \nr00071[31] [18] : \nr00071[30] [18];
  assign nw03861 = nr00001[1] ? nw03860 : nw03859;
  assign nw03862 = nr00001[2] ? nw03861 : nw03858;
  assign nw03863 = nr00001[3] ? nw03862 : nw03855;
  assign nw00179 = nr00001[4] ? nw03863 : nw03848;
  assign nw00326 = nw03323 ? \nr00067 [18] : nw00179;
  assign nw03864 = nr00001[0] ? \nr00071[1] [19] : \nr00071[0] [19];
  assign nw03865 = nr00001[0] ? \nr00071[3] [19] : \nr00071[2] [19];
  assign nw03866 = nr00001[1] ? nw03865 : nw03864;
  assign nw03867 = nr00001[0] ? \nr00071[5] [19] : \nr00071[4] [19];
  assign nw03868 = nr00001[0] ? \nr00071[7] [19] : \nr00071[6] [19];
  assign nw03869 = nr00001[1] ? nw03868 : nw03867;
  assign nw03870 = nr00001[2] ? nw03869 : nw03866;
  assign nw03871 = nr00001[0] ? \nr00071[9] [19] : \nr00071[8] [19];
  assign nw03872 = nr00001[0] ? \nr00071[11] [19] : \nr00071[10] [19];
  assign nw03873 = nr00001[1] ? nw03872 : nw03871;
  assign nw03874 = nr00001[0] ? \nr00071[13] [19] : \nr00071[12] [19];
  assign nw03875 = nr00001[0] ? \nr00071[15] [19] : \nr00071[14] [19];
  assign nw03876 = nr00001[1] ? nw03875 : nw03874;
  assign nw03877 = nr00001[2] ? nw03876 : nw03873;
  assign nw03878 = nr00001[3] ? nw03877 : nw03870;
  assign nw03879 = nr00001[0] ? \nr00071[17] [19] : \nr00071[16] [19];
  assign nw03880 = nr00001[0] ? \nr00071[19] [19] : \nr00071[18] [19];
  assign nw03881 = nr00001[1] ? nw03880 : nw03879;
  assign nw03882 = nr00001[0] ? \nr00071[21] [19] : \nr00071[20] [19];
  assign nw03883 = nr00001[0] ? \nr00071[23] [19] : \nr00071[22] [19];
  assign nw03884 = nr00001[1] ? nw03883 : nw03882;
  assign nw03885 = nr00001[2] ? nw03884 : nw03881;
  assign nw03886 = nr00001[0] ? \nr00071[25] [19] : \nr00071[24] [19];
  assign nw03887 = nr00001[0] ? \nr00071[27] [19] : \nr00071[26] [19];
  assign nw03888 = nr00001[1] ? nw03887 : nw03886;
  assign nw03889 = nr00001[0] ? \nr00071[29] [19] : \nr00071[28] [19];
  assign nw03890 = nr00001[0] ? \nr00071[31] [19] : \nr00071[30] [19];
  assign nw03891 = nr00001[1] ? nw03890 : nw03889;
  assign nw03892 = nr00001[2] ? nw03891 : nw03888;
  assign nw03893 = nr00001[3] ? nw03892 : nw03885;
  assign nw00180 = nr00001[4] ? nw03893 : nw03878;
  assign nw00327 = nw03323 ? \nr00067 [19] : nw00180;
  assign nw03894 = nr00001[0] ? \nr00071[1] [20] : \nr00071[0] [20];
  assign nw03895 = nr00001[0] ? \nr00071[3] [20] : \nr00071[2] [20];
  assign nw03896 = nr00001[1] ? nw03895 : nw03894;
  assign nw03897 = nr00001[0] ? \nr00071[5] [20] : \nr00071[4] [20];
  assign nw03898 = nr00001[0] ? \nr00071[7] [20] : \nr00071[6] [20];
  assign nw03899 = nr00001[1] ? nw03898 : nw03897;
  assign nw03900 = nr00001[2] ? nw03899 : nw03896;
  assign nw03901 = nr00001[0] ? \nr00071[9] [20] : \nr00071[8] [20];
  assign nw03902 = nr00001[0] ? \nr00071[11] [20] : \nr00071[10] [20];
  assign nw03903 = nr00001[1] ? nw03902 : nw03901;
  assign nw03904 = nr00001[0] ? \nr00071[13] [20] : \nr00071[12] [20];
  assign nw03905 = nr00001[0] ? \nr00071[15] [20] : \nr00071[14] [20];
  assign nw03906 = nr00001[1] ? nw03905 : nw03904;
  assign nw03907 = nr00001[2] ? nw03906 : nw03903;
  assign nw03908 = nr00001[3] ? nw03907 : nw03900;
  assign nw03909 = nr00001[0] ? \nr00071[17] [20] : \nr00071[16] [20];
  assign nw03910 = nr00001[0] ? \nr00071[19] [20] : \nr00071[18] [20];
  assign nw03911 = nr00001[1] ? nw03910 : nw03909;
  assign nw03912 = nr00001[0] ? \nr00071[21] [20] : \nr00071[20] [20];
  assign nw03913 = nr00001[0] ? \nr00071[23] [20] : \nr00071[22] [20];
  assign nw03914 = nr00001[1] ? nw03913 : nw03912;
  assign nw03915 = nr00001[2] ? nw03914 : nw03911;
  assign nw03916 = nr00001[0] ? \nr00071[25] [20] : \nr00071[24] [20];
  assign nw03917 = nr00001[0] ? \nr00071[27] [20] : \nr00071[26] [20];
  assign nw03918 = nr00001[1] ? nw03917 : nw03916;
  assign nw03919 = nr00001[0] ? \nr00071[29] [20] : \nr00071[28] [20];
  assign nw03920 = nr00001[0] ? \nr00071[31] [20] : \nr00071[30] [20];
  assign nw03921 = nr00001[1] ? nw03920 : nw03919;
  assign nw03922 = nr00001[2] ? nw03921 : nw03918;
  assign nw03923 = nr00001[3] ? nw03922 : nw03915;
  assign nw00182 = nr00001[4] ? nw03923 : nw03908;
  assign nw00329 = nw03323 ? \nr00067 [20] : nw00182;
  assign nw03924 = nr00001[0] ? \nr00071[1] [21] : \nr00071[0] [21];
  assign nw03925 = nr00001[0] ? \nr00071[3] [21] : \nr00071[2] [21];
  assign nw03926 = nr00001[1] ? nw03925 : nw03924;
  assign nw03927 = nr00001[0] ? \nr00071[5] [21] : \nr00071[4] [21];
  assign nw03928 = nr00001[0] ? \nr00071[7] [21] : \nr00071[6] [21];
  assign nw03929 = nr00001[1] ? nw03928 : nw03927;
  assign nw03930 = nr00001[2] ? nw03929 : nw03926;
  assign nw03931 = nr00001[0] ? \nr00071[9] [21] : \nr00071[8] [21];
  assign nw03932 = nr00001[0] ? \nr00071[11] [21] : \nr00071[10] [21];
  assign nw03933 = nr00001[1] ? nw03932 : nw03931;
  assign nw03934 = nr00001[0] ? \nr00071[13] [21] : \nr00071[12] [21];
  assign nw03935 = nr00001[0] ? \nr00071[15] [21] : \nr00071[14] [21];
  assign nw03936 = nr00001[1] ? nw03935 : nw03934;
  assign nw03937 = nr00001[2] ? nw03936 : nw03933;
  assign nw03938 = nr00001[3] ? nw03937 : nw03930;
  assign nw03939 = nr00001[0] ? \nr00071[17] [21] : \nr00071[16] [21];
  assign nw03940 = nr00001[0] ? \nr00071[19] [21] : \nr00071[18] [21];
  assign nw03941 = nr00001[1] ? nw03940 : nw03939;
  assign nw03942 = nr00001[0] ? \nr00071[21] [21] : \nr00071[20] [21];
  assign nw03943 = nr00001[0] ? \nr00071[23] [21] : \nr00071[22] [21];
  assign nw03944 = nr00001[1] ? nw03943 : nw03942;
  assign nw03945 = nr00001[2] ? nw03944 : nw03941;
  assign nw03946 = nr00001[0] ? \nr00071[25] [21] : \nr00071[24] [21];
  assign nw03947 = nr00001[0] ? \nr00071[27] [21] : \nr00071[26] [21];
  assign nw03948 = nr00001[1] ? nw03947 : nw03946;
  assign nw03949 = nr00001[0] ? \nr00071[29] [21] : \nr00071[28] [21];
  assign nw03950 = nr00001[0] ? \nr00071[31] [21] : \nr00071[30] [21];
  assign nw03951 = nr00001[1] ? nw03950 : nw03949;
  assign nw03952 = nr00001[2] ? nw03951 : nw03948;
  assign nw03953 = nr00001[3] ? nw03952 : nw03945;
  assign nw00183 = nr00001[4] ? nw03953 : nw03938;
  assign nw00330 = nw03323 ? \nr00067 [21] : nw00183;
  assign nw03954 = nr00001[0] ? \nr00071[1] [22] : \nr00071[0] [22];
  assign nw03955 = nr00001[0] ? \nr00071[3] [22] : \nr00071[2] [22];
  assign nw03956 = nr00001[1] ? nw03955 : nw03954;
  assign nw03957 = nr00001[0] ? \nr00071[5] [22] : \nr00071[4] [22];
  assign nw03958 = nr00001[0] ? \nr00071[7] [22] : \nr00071[6] [22];
  assign nw03959 = nr00001[1] ? nw03958 : nw03957;
  assign nw03960 = nr00001[2] ? nw03959 : nw03956;
  assign nw03961 = nr00001[0] ? \nr00071[9] [22] : \nr00071[8] [22];
  assign nw03962 = nr00001[0] ? \nr00071[11] [22] : \nr00071[10] [22];
  assign nw03963 = nr00001[1] ? nw03962 : nw03961;
  assign nw03964 = nr00001[0] ? \nr00071[13] [22] : \nr00071[12] [22];
  assign nw03965 = nr00001[0] ? \nr00071[15] [22] : \nr00071[14] [22];
  assign nw03966 = nr00001[1] ? nw03965 : nw03964;
  assign nw03967 = nr00001[2] ? nw03966 : nw03963;
  assign nw03968 = nr00001[3] ? nw03967 : nw03960;
  assign nw03969 = nr00001[0] ? \nr00071[17] [22] : \nr00071[16] [22];
  assign nw03970 = nr00001[0] ? \nr00071[19] [22] : \nr00071[18] [22];
  assign nw03971 = nr00001[1] ? nw03970 : nw03969;
  assign nw03972 = nr00001[0] ? \nr00071[21] [22] : \nr00071[20] [22];
  assign nw03973 = nr00001[0] ? \nr00071[23] [22] : \nr00071[22] [22];
  assign nw03974 = nr00001[1] ? nw03973 : nw03972;
  assign nw03975 = nr00001[2] ? nw03974 : nw03971;
  assign nw03976 = nr00001[0] ? \nr00071[25] [22] : \nr00071[24] [22];
  assign nw03977 = nr00001[0] ? \nr00071[27] [22] : \nr00071[26] [22];
  assign nw03978 = nr00001[1] ? nw03977 : nw03976;
  assign nw03979 = nr00001[0] ? \nr00071[29] [22] : \nr00071[28] [22];
  assign nw03980 = nr00001[0] ? \nr00071[31] [22] : \nr00071[30] [22];
  assign nw03981 = nr00001[1] ? nw03980 : nw03979;
  assign nw03982 = nr00001[2] ? nw03981 : nw03978;
  assign nw03983 = nr00001[3] ? nw03982 : nw03975;
  assign nw00184 = nr00001[4] ? nw03983 : nw03968;
  assign nw00331 = nw03323 ? \nr00067 [22] : nw00184;
  assign nw03984 = nr00001[0] ? \nr00071[1] [23] : \nr00071[0] [23];
  assign nw03985 = nr00001[0] ? \nr00071[3] [23] : \nr00071[2] [23];
  assign nw03986 = nr00001[1] ? nw03985 : nw03984;
  assign nw03987 = nr00001[0] ? \nr00071[5] [23] : \nr00071[4] [23];
  assign nw03988 = nr00001[0] ? \nr00071[7] [23] : \nr00071[6] [23];
  assign nw03989 = nr00001[1] ? nw03988 : nw03987;
  assign nw03990 = nr00001[2] ? nw03989 : nw03986;
  assign nw03991 = nr00001[0] ? \nr00071[9] [23] : \nr00071[8] [23];
  assign nw03992 = nr00001[0] ? \nr00071[11] [23] : \nr00071[10] [23];
  assign nw03993 = nr00001[1] ? nw03992 : nw03991;
  assign nw03994 = nr00001[0] ? \nr00071[13] [23] : \nr00071[12] [23];
  assign nw03995 = nr00001[0] ? \nr00071[15] [23] : \nr00071[14] [23];
  assign nw03996 = nr00001[1] ? nw03995 : nw03994;
  assign nw03997 = nr00001[2] ? nw03996 : nw03993;
  assign nw03998 = nr00001[3] ? nw03997 : nw03990;
  assign nw03999 = nr00001[0] ? \nr00071[17] [23] : \nr00071[16] [23];
  assign nw04000 = nr00001[0] ? \nr00071[19] [23] : \nr00071[18] [23];
  assign nw04001 = nr00001[1] ? nw04000 : nw03999;
  assign nw04002 = nr00001[0] ? \nr00071[21] [23] : \nr00071[20] [23];
  assign nw04003 = nr00001[0] ? \nr00071[23] [23] : \nr00071[22] [23];
  assign nw04004 = nr00001[1] ? nw04003 : nw04002;
  assign nw04005 = nr00001[2] ? nw04004 : nw04001;
  assign nw04006 = nr00001[0] ? \nr00071[25] [23] : \nr00071[24] [23];
  assign nw04007 = nr00001[0] ? \nr00071[27] [23] : \nr00071[26] [23];
  assign nw04008 = nr00001[1] ? nw04007 : nw04006;
  assign nw04009 = nr00001[0] ? \nr00071[29] [23] : \nr00071[28] [23];
  assign nw04010 = nr00001[0] ? \nr00071[31] [23] : \nr00071[30] [23];
  assign nw04011 = nr00001[1] ? nw04010 : nw04009;
  assign nw04012 = nr00001[2] ? nw04011 : nw04008;
  assign nw04013 = nr00001[3] ? nw04012 : nw04005;
  assign nw00185 = nr00001[4] ? nw04013 : nw03998;
  assign nw00332 = nw03323 ? \nr00067 [23] : nw00185;
  assign nw04014 = nr00001[0] ? \nr00071[1] [24] : \nr00071[0] [24];
  assign nw04015 = nr00001[0] ? \nr00071[3] [24] : \nr00071[2] [24];
  assign nw04016 = nr00001[1] ? nw04015 : nw04014;
  assign nw04017 = nr00001[0] ? \nr00071[5] [24] : \nr00071[4] [24];
  assign nw04018 = nr00001[0] ? \nr00071[7] [24] : \nr00071[6] [24];
  assign nw04019 = nr00001[1] ? nw04018 : nw04017;
  assign nw04020 = nr00001[2] ? nw04019 : nw04016;
  assign nw04021 = nr00001[0] ? \nr00071[9] [24] : \nr00071[8] [24];
  assign nw04022 = nr00001[0] ? \nr00071[11] [24] : \nr00071[10] [24];
  assign nw04023 = nr00001[1] ? nw04022 : nw04021;
  assign nw04024 = nr00001[0] ? \nr00071[13] [24] : \nr00071[12] [24];
  assign nw04025 = nr00001[0] ? \nr00071[15] [24] : \nr00071[14] [24];
  assign nw04026 = nr00001[1] ? nw04025 : nw04024;
  assign nw04027 = nr00001[2] ? nw04026 : nw04023;
  assign nw04028 = nr00001[3] ? nw04027 : nw04020;
  assign nw04029 = nr00001[0] ? \nr00071[17] [24] : \nr00071[16] [24];
  assign nw04030 = nr00001[0] ? \nr00071[19] [24] : \nr00071[18] [24];
  assign nw04031 = nr00001[1] ? nw04030 : nw04029;
  assign nw04032 = nr00001[0] ? \nr00071[21] [24] : \nr00071[20] [24];
  assign nw04033 = nr00001[0] ? \nr00071[23] [24] : \nr00071[22] [24];
  assign nw04034 = nr00001[1] ? nw04033 : nw04032;
  assign nw04035 = nr00001[2] ? nw04034 : nw04031;
  assign nw04036 = nr00001[0] ? \nr00071[25] [24] : \nr00071[24] [24];
  assign nw04037 = nr00001[0] ? \nr00071[27] [24] : \nr00071[26] [24];
  assign nw04038 = nr00001[1] ? nw04037 : nw04036;
  assign nw04039 = nr00001[0] ? \nr00071[29] [24] : \nr00071[28] [24];
  assign nw04040 = nr00001[0] ? \nr00071[31] [24] : \nr00071[30] [24];
  assign nw04041 = nr00001[1] ? nw04040 : nw04039;
  assign nw04042 = nr00001[2] ? nw04041 : nw04038;
  assign nw04043 = nr00001[3] ? nw04042 : nw04035;
  assign nw00186 = nr00001[4] ? nw04043 : nw04028;
  assign nw00333 = nw03323 ? \nr00067 [24] : nw00186;
  assign nw04044 = nr00001[0] ? \nr00071[1] [25] : \nr00071[0] [25];
  assign nw04045 = nr00001[0] ? \nr00071[3] [25] : \nr00071[2] [25];
  assign nw04046 = nr00001[1] ? nw04045 : nw04044;
  assign nw04047 = nr00001[0] ? \nr00071[5] [25] : \nr00071[4] [25];
  assign nw04048 = nr00001[0] ? \nr00071[7] [25] : \nr00071[6] [25];
  assign nw04049 = nr00001[1] ? nw04048 : nw04047;
  assign nw04050 = nr00001[2] ? nw04049 : nw04046;
  assign nw04051 = nr00001[0] ? \nr00071[9] [25] : \nr00071[8] [25];
  assign nw04052 = nr00001[0] ? \nr00071[11] [25] : \nr00071[10] [25];
  assign nw04053 = nr00001[1] ? nw04052 : nw04051;
  assign nw04054 = nr00001[0] ? \nr00071[13] [25] : \nr00071[12] [25];
  assign nw04055 = nr00001[0] ? \nr00071[15] [25] : \nr00071[14] [25];
  assign nw04056 = nr00001[1] ? nw04055 : nw04054;
  assign nw04057 = nr00001[2] ? nw04056 : nw04053;
  assign nw04058 = nr00001[3] ? nw04057 : nw04050;
  assign nw04059 = nr00001[0] ? \nr00071[17] [25] : \nr00071[16] [25];
  assign nw04060 = nr00001[0] ? \nr00071[19] [25] : \nr00071[18] [25];
  assign nw04061 = nr00001[1] ? nw04060 : nw04059;
  assign nw04062 = nr00001[0] ? \nr00071[21] [25] : \nr00071[20] [25];
  assign nw04063 = nr00001[0] ? \nr00071[23] [25] : \nr00071[22] [25];
  assign nw04064 = nr00001[1] ? nw04063 : nw04062;
  assign nw04065 = nr00001[2] ? nw04064 : nw04061;
  assign nw04066 = nr00001[0] ? \nr00071[25] [25] : \nr00071[24] [25];
  assign nw04067 = nr00001[0] ? \nr00071[27] [25] : \nr00071[26] [25];
  assign nw04068 = nr00001[1] ? nw04067 : nw04066;
  assign nw04069 = nr00001[0] ? \nr00071[29] [25] : \nr00071[28] [25];
  assign nw04070 = nr00001[0] ? \nr00071[31] [25] : \nr00071[30] [25];
  assign nw04071 = nr00001[1] ? nw04070 : nw04069;
  assign nw04072 = nr00001[2] ? nw04071 : nw04068;
  assign nw04073 = nr00001[3] ? nw04072 : nw04065;
  assign nw00187 = nr00001[4] ? nw04073 : nw04058;
  assign nw00334 = nw03323 ? \nr00067 [25] : nw00187;
  assign nw04074 = nr00001[0] ? \nr00071[1] [26] : \nr00071[0] [26];
  assign nw04075 = nr00001[0] ? \nr00071[3] [26] : \nr00071[2] [26];
  assign nw04076 = nr00001[1] ? nw04075 : nw04074;
  assign nw04077 = nr00001[0] ? \nr00071[5] [26] : \nr00071[4] [26];
  assign nw04078 = nr00001[0] ? \nr00071[7] [26] : \nr00071[6] [26];
  assign nw04079 = nr00001[1] ? nw04078 : nw04077;
  assign nw04080 = nr00001[2] ? nw04079 : nw04076;
  assign nw04081 = nr00001[0] ? \nr00071[9] [26] : \nr00071[8] [26];
  assign nw04082 = nr00001[0] ? \nr00071[11] [26] : \nr00071[10] [26];
  assign nw04083 = nr00001[1] ? nw04082 : nw04081;
  assign nw04084 = nr00001[0] ? \nr00071[13] [26] : \nr00071[12] [26];
  assign nw04085 = nr00001[0] ? \nr00071[15] [26] : \nr00071[14] [26];
  assign nw04086 = nr00001[1] ? nw04085 : nw04084;
  assign nw04087 = nr00001[2] ? nw04086 : nw04083;
  assign nw04088 = nr00001[3] ? nw04087 : nw04080;
  assign nw04089 = nr00001[0] ? \nr00071[17] [26] : \nr00071[16] [26];
  assign nw04090 = nr00001[0] ? \nr00071[19] [26] : \nr00071[18] [26];
  assign nw04091 = nr00001[1] ? nw04090 : nw04089;
  assign nw04092 = nr00001[0] ? \nr00071[21] [26] : \nr00071[20] [26];
  assign nw04093 = nr00001[0] ? \nr00071[23] [26] : \nr00071[22] [26];
  assign nw04094 = nr00001[1] ? nw04093 : nw04092;
  assign nw04095 = nr00001[2] ? nw04094 : nw04091;
  assign nw04096 = nr00001[0] ? \nr00071[25] [26] : \nr00071[24] [26];
  assign nw04097 = nr00001[0] ? \nr00071[27] [26] : \nr00071[26] [26];
  assign nw04098 = nr00001[1] ? nw04097 : nw04096;
  assign nw04099 = nr00001[0] ? \nr00071[29] [26] : \nr00071[28] [26];
  assign nw04100 = nr00001[0] ? \nr00071[31] [26] : \nr00071[30] [26];
  assign nw04101 = nr00001[1] ? nw04100 : nw04099;
  assign nw04102 = nr00001[2] ? nw04101 : nw04098;
  assign nw04103 = nr00001[3] ? nw04102 : nw04095;
  assign nw00188 = nr00001[4] ? nw04103 : nw04088;
  assign nw00335 = nw03323 ? \nr00067 [26] : nw00188;
  assign nw04104 = nr00001[0] ? \nr00071[1] [27] : \nr00071[0] [27];
  assign nw04105 = nr00001[0] ? \nr00071[3] [27] : \nr00071[2] [27];
  assign nw04106 = nr00001[1] ? nw04105 : nw04104;
  assign nw04107 = nr00001[0] ? \nr00071[5] [27] : \nr00071[4] [27];
  assign nw04108 = nr00001[0] ? \nr00071[7] [27] : \nr00071[6] [27];
  assign nw04109 = nr00001[1] ? nw04108 : nw04107;
  assign nw04110 = nr00001[2] ? nw04109 : nw04106;
  assign nw04111 = nr00001[0] ? \nr00071[9] [27] : \nr00071[8] [27];
  assign nw04112 = nr00001[0] ? \nr00071[11] [27] : \nr00071[10] [27];
  assign nw04113 = nr00001[1] ? nw04112 : nw04111;
  assign nw04114 = nr00001[0] ? \nr00071[13] [27] : \nr00071[12] [27];
  assign nw04115 = nr00001[0] ? \nr00071[15] [27] : \nr00071[14] [27];
  assign nw04116 = nr00001[1] ? nw04115 : nw04114;
  assign nw04117 = nr00001[2] ? nw04116 : nw04113;
  assign nw04118 = nr00001[3] ? nw04117 : nw04110;
  assign nw04119 = nr00001[0] ? \nr00071[17] [27] : \nr00071[16] [27];
  assign nw04120 = nr00001[0] ? \nr00071[19] [27] : \nr00071[18] [27];
  assign nw04121 = nr00001[1] ? nw04120 : nw04119;
  assign nw04122 = nr00001[0] ? \nr00071[21] [27] : \nr00071[20] [27];
  assign nw04123 = nr00001[0] ? \nr00071[23] [27] : \nr00071[22] [27];
  assign nw04124 = nr00001[1] ? nw04123 : nw04122;
  assign nw04125 = nr00001[2] ? nw04124 : nw04121;
  assign nw04126 = nr00001[0] ? \nr00071[25] [27] : \nr00071[24] [27];
  assign nw04127 = nr00001[0] ? \nr00071[27] [27] : \nr00071[26] [27];
  assign nw04128 = nr00001[1] ? nw04127 : nw04126;
  assign nw04129 = nr00001[0] ? \nr00071[29] [27] : \nr00071[28] [27];
  assign nw04130 = nr00001[0] ? \nr00071[31] [27] : \nr00071[30] [27];
  assign nw04131 = nr00001[1] ? nw04130 : nw04129;
  assign nw04132 = nr00001[2] ? nw04131 : nw04128;
  assign nw04133 = nr00001[3] ? nw04132 : nw04125;
  assign nw00189 = nr00001[4] ? nw04133 : nw04118;
  assign nw00336 = nw03323 ? \nr00067 [27] : nw00189;
  assign nw04134 = nr00001[0] ? \nr00071[1] [28] : \nr00071[0] [28];
  assign nw04135 = nr00001[0] ? \nr00071[3] [28] : \nr00071[2] [28];
  assign nw04136 = nr00001[1] ? nw04135 : nw04134;
  assign nw04137 = nr00001[0] ? \nr00071[5] [28] : \nr00071[4] [28];
  assign nw04138 = nr00001[0] ? \nr00071[7] [28] : \nr00071[6] [28];
  assign nw04139 = nr00001[1] ? nw04138 : nw04137;
  assign nw04140 = nr00001[2] ? nw04139 : nw04136;
  assign nw04141 = nr00001[0] ? \nr00071[9] [28] : \nr00071[8] [28];
  assign nw04142 = nr00001[0] ? \nr00071[11] [28] : \nr00071[10] [28];
  assign nw04143 = nr00001[1] ? nw04142 : nw04141;
  assign nw04144 = nr00001[0] ? \nr00071[13] [28] : \nr00071[12] [28];
  assign nw04145 = nr00001[0] ? \nr00071[15] [28] : \nr00071[14] [28];
  assign nw04146 = nr00001[1] ? nw04145 : nw04144;
  assign nw04147 = nr00001[2] ? nw04146 : nw04143;
  assign nw04148 = nr00001[3] ? nw04147 : nw04140;
  assign nw04149 = nr00001[0] ? \nr00071[17] [28] : \nr00071[16] [28];
  assign nw04150 = nr00001[0] ? \nr00071[19] [28] : \nr00071[18] [28];
  assign nw04151 = nr00001[1] ? nw04150 : nw04149;
  assign nw04152 = nr00001[0] ? \nr00071[21] [28] : \nr00071[20] [28];
  assign nw04153 = nr00001[0] ? \nr00071[23] [28] : \nr00071[22] [28];
  assign nw04154 = nr00001[1] ? nw04153 : nw04152;
  assign nw04155 = nr00001[2] ? nw04154 : nw04151;
  assign nw04156 = nr00001[0] ? \nr00071[25] [28] : \nr00071[24] [28];
  assign nw04157 = nr00001[0] ? \nr00071[27] [28] : \nr00071[26] [28];
  assign nw04158 = nr00001[1] ? nw04157 : nw04156;
  assign nw04159 = nr00001[0] ? \nr00071[29] [28] : \nr00071[28] [28];
  assign nw04160 = nr00001[0] ? \nr00071[31] [28] : \nr00071[30] [28];
  assign nw04161 = nr00001[1] ? nw04160 : nw04159;
  assign nw04162 = nr00001[2] ? nw04161 : nw04158;
  assign nw04163 = nr00001[3] ? nw04162 : nw04155;
  assign nw00190 = nr00001[4] ? nw04163 : nw04148;
  assign nw00337 = nw03323 ? \nr00067 [28] : nw00190;
  assign nw04164 = nr00001[0] ? \nr00071[1] [29] : \nr00071[0] [29];
  assign nw04165 = nr00001[0] ? \nr00071[3] [29] : \nr00071[2] [29];
  assign nw04166 = nr00001[1] ? nw04165 : nw04164;
  assign nw04167 = nr00001[0] ? \nr00071[5] [29] : \nr00071[4] [29];
  assign nw04168 = nr00001[0] ? \nr00071[7] [29] : \nr00071[6] [29];
  assign nw04169 = nr00001[1] ? nw04168 : nw04167;
  assign nw04170 = nr00001[2] ? nw04169 : nw04166;
  assign nw04171 = nr00001[0] ? \nr00071[9] [29] : \nr00071[8] [29];
  assign nw04172 = nr00001[0] ? \nr00071[11] [29] : \nr00071[10] [29];
  assign nw04173 = nr00001[1] ? nw04172 : nw04171;
  assign nw04174 = nr00001[0] ? \nr00071[13] [29] : \nr00071[12] [29];
  assign nw04175 = nr00001[0] ? \nr00071[15] [29] : \nr00071[14] [29];
  assign nw04176 = nr00001[1] ? nw04175 : nw04174;
  assign nw04177 = nr00001[2] ? nw04176 : nw04173;
  assign nw04178 = nr00001[3] ? nw04177 : nw04170;
  assign nw04179 = nr00001[0] ? \nr00071[17] [29] : \nr00071[16] [29];
  assign nw04180 = nr00001[0] ? \nr00071[19] [29] : \nr00071[18] [29];
  assign nw04181 = nr00001[1] ? nw04180 : nw04179;
  assign nw04182 = nr00001[0] ? \nr00071[21] [29] : \nr00071[20] [29];
  assign nw04183 = nr00001[0] ? \nr00071[23] [29] : \nr00071[22] [29];
  assign nw04184 = nr00001[1] ? nw04183 : nw04182;
  assign nw04185 = nr00001[2] ? nw04184 : nw04181;
  assign nw04186 = nr00001[0] ? \nr00071[25] [29] : \nr00071[24] [29];
  assign nw04187 = nr00001[0] ? \nr00071[27] [29] : \nr00071[26] [29];
  assign nw04188 = nr00001[1] ? nw04187 : nw04186;
  assign nw04189 = nr00001[0] ? \nr00071[29] [29] : \nr00071[28] [29];
  assign nw04190 = nr00001[0] ? \nr00071[31] [29] : \nr00071[30] [29];
  assign nw04191 = nr00001[1] ? nw04190 : nw04189;
  assign nw04192 = nr00001[2] ? nw04191 : nw04188;
  assign nw04193 = nr00001[3] ? nw04192 : nw04185;
  assign nw00191 = nr00001[4] ? nw04193 : nw04178;
  assign nw00338 = nw03323 ? \nr00067 [29] : nw00191;
  assign nw04194 = nr00001[0] ? \nr00071[1] [30] : \nr00071[0] [30];
  assign nw04195 = nr00001[0] ? \nr00071[3] [30] : \nr00071[2] [30];
  assign nw04196 = nr00001[1] ? nw04195 : nw04194;
  assign nw04197 = nr00001[0] ? \nr00071[5] [30] : \nr00071[4] [30];
  assign nw04198 = nr00001[0] ? \nr00071[7] [30] : \nr00071[6] [30];
  assign nw04199 = nr00001[1] ? nw04198 : nw04197;
  assign nw04200 = nr00001[2] ? nw04199 : nw04196;
  assign nw04201 = nr00001[0] ? \nr00071[9] [30] : \nr00071[8] [30];
  assign nw04202 = nr00001[0] ? \nr00071[11] [30] : \nr00071[10] [30];
  assign nw04203 = nr00001[1] ? nw04202 : nw04201;
  assign nw04204 = nr00001[0] ? \nr00071[13] [30] : \nr00071[12] [30];
  assign nw04205 = nr00001[0] ? \nr00071[15] [30] : \nr00071[14] [30];
  assign nw04206 = nr00001[1] ? nw04205 : nw04204;
  assign nw04207 = nr00001[2] ? nw04206 : nw04203;
  assign nw04208 = nr00001[3] ? nw04207 : nw04200;
  assign nw04209 = nr00001[0] ? \nr00071[17] [30] : \nr00071[16] [30];
  assign nw04210 = nr00001[0] ? \nr00071[19] [30] : \nr00071[18] [30];
  assign nw04211 = nr00001[1] ? nw04210 : nw04209;
  assign nw04212 = nr00001[0] ? \nr00071[21] [30] : \nr00071[20] [30];
  assign nw04213 = nr00001[0] ? \nr00071[23] [30] : \nr00071[22] [30];
  assign nw04214 = nr00001[1] ? nw04213 : nw04212;
  assign nw04215 = nr00001[2] ? nw04214 : nw04211;
  assign nw04216 = nr00001[0] ? \nr00071[25] [30] : \nr00071[24] [30];
  assign nw04217 = nr00001[0] ? \nr00071[27] [30] : \nr00071[26] [30];
  assign nw04218 = nr00001[1] ? nw04217 : nw04216;
  assign nw04219 = nr00001[0] ? \nr00071[29] [30] : \nr00071[28] [30];
  assign nw04220 = nr00001[0] ? \nr00071[31] [30] : \nr00071[30] [30];
  assign nw04221 = nr00001[1] ? nw04220 : nw04219;
  assign nw04222 = nr00001[2] ? nw04221 : nw04218;
  assign nw04223 = nr00001[3] ? nw04222 : nw04215;
  assign nw00193 = nr00001[4] ? nw04223 : nw04208;
  assign nw00340 = nw03323 ? \nr00067 [30] : nw00193;
  assign nw04224 = nr00001[0] ? \nr00071[1] [31] : \nr00071[0] [31];
  assign nw04225 = nr00001[0] ? \nr00071[3] [31] : \nr00071[2] [31];
  assign nw04226 = nr00001[1] ? nw04225 : nw04224;
  assign nw04227 = nr00001[0] ? \nr00071[5] [31] : \nr00071[4] [31];
  assign nw04228 = nr00001[0] ? \nr00071[7] [31] : \nr00071[6] [31];
  assign nw04229 = nr00001[1] ? nw04228 : nw04227;
  assign nw04230 = nr00001[2] ? nw04229 : nw04226;
  assign nw04231 = nr00001[0] ? \nr00071[9] [31] : \nr00071[8] [31];
  assign nw04232 = nr00001[0] ? \nr00071[11] [31] : \nr00071[10] [31];
  assign nw04233 = nr00001[1] ? nw04232 : nw04231;
  assign nw04234 = nr00001[0] ? \nr00071[13] [31] : \nr00071[12] [31];
  assign nw04235 = nr00001[0] ? \nr00071[15] [31] : \nr00071[14] [31];
  assign nw04236 = nr00001[1] ? nw04235 : nw04234;
  assign nw04237 = nr00001[2] ? nw04236 : nw04233;
  assign nw04238 = nr00001[3] ? nw04237 : nw04230;
  assign nw04239 = nr00001[0] ? \nr00071[17] [31] : \nr00071[16] [31];
  assign nw04240 = nr00001[0] ? \nr00071[19] [31] : \nr00071[18] [31];
  assign nw04241 = nr00001[1] ? nw04240 : nw04239;
  assign nw04242 = nr00001[0] ? \nr00071[21] [31] : \nr00071[20] [31];
  assign nw04243 = nr00001[0] ? \nr00071[23] [31] : \nr00071[22] [31];
  assign nw04244 = nr00001[1] ? nw04243 : nw04242;
  assign nw04245 = nr00001[2] ? nw04244 : nw04241;
  assign nw04246 = nr00001[0] ? \nr00071[25] [31] : \nr00071[24] [31];
  assign nw04247 = nr00001[0] ? \nr00071[27] [31] : \nr00071[26] [31];
  assign nw04248 = nr00001[1] ? nw04247 : nw04246;
  assign nw04249 = nr00001[0] ? \nr00071[29] [31] : \nr00071[28] [31];
  assign nw04250 = nr00001[0] ? \nr00071[31] [31] : \nr00071[30] [31];
  assign nw04251 = nr00001[1] ? nw04250 : nw04249;
  assign nw04252 = nr00001[2] ? nw04251 : nw04248;
  assign nw04253 = nr00001[3] ? nw04252 : nw04245;
  assign nw00194 = nr00001[4] ? nw04253 : nw04238;
  assign nw00341 = nw03323 ? \nr00067 [31] : nw00194;
  assign nw04254 = \nr00050I  | \nr00058I ;
  assign \nw05426  = nw04254 | \nr00056I ;
  assign nw04255 = \nr00027  | \nr00015 ;
  assign nw04256 = nw04255 | \nr00052 ;
  assign nw04257 = nw04256 | \nr00052U ;
  assign nw04258 = nw04257 | \nr00061 ;
  assign nw04259 = ~(nw04258 | \nr00046 );
  assign nw04260 = nw04259 & ~(\nr00028 );
  assign nw04261 = \nr00050  | \nr00058 ;
  assign nw04262 = nw04261 | \nr00056 ;
  assign nw04263 = nw04260 & ~(nw04262);
  assign nw04264 = nw04263 ? \nr00026 [0] : nw00202;
  assign nw00097 = \nw05426  ? \nr00070 [0] : nw04264;
  assign nw04265 = nw04263 ? \nr00026 [1] : nw00213;
  assign nw00098 = \nw05426  ? \nr00070 [1] : nw04265;
  assign nw04266 = nw04263 ? \nr00026 [2] : nw00224;
  assign nw00099 = \nw05426  ? \nr00070 [2] : nw04266;
  assign nw04267 = nw04263 ? \nr00026 [3] : nw00227;
  assign nw00100 = \nw05426  ? \nr00070 [3] : nw04267;
  assign nw04268 = nw04263 ? \nr00026 [4] : nw00228;
  assign nw00101 = \nw05426  ? \nr00070 [4] : nw04268;
  assign nw00312 = nw04263 ? \nr00026 [5] : nw00229;
  assign nw00313 = nw04263 ? \nr00026 [6] : nw00230;
  assign nw00314 = nw04263 ? \nr00026 [7] : nw00231;
  assign nw00315 = nw04263 ? \nr00026 [8] : nw00232;
  assign nw00316 = nw04263 ? \nr00026 [9] : nw00233;
  assign nw00290 = nw04263 ? \nr00026 [10] : nw00203;
  assign nw00291 = nw04263 ? \nr00026 [11] : nw00204;
  assign nw00292 = nw04263 ? \nr00026 [12] : nw00205;
  assign nw00293 = nw04263 ? \nr00026 [13] : nw00206;
  assign nw00294 = nw04263 ? \nr00026 [14] : nw00207;
  assign nw00295 = nw04263 ? \nr00026 [15] : nw00208;
  assign nw00296 = nw04263 ? \nr00026 [16] : nw00209;
  assign nw00297 = nw04263 ? \nr00026 [17] : nw00210;
  assign nw00298 = nw04263 ? \nr00026 [18] : nw00211;
  assign nw00299 = nw04263 ? \nr00026 [19] : nw00212;
  assign nw00300 = nw04263 ? \nr00026 [20] : nw00214;
  assign nw00301 = nw04263 ? \nr00026 [21] : nw00215;
  assign nw00302 = nw04263 ? \nr00026 [22] : nw00216;
  assign nw00303 = nw04263 ? \nr00026 [23] : nw00217;
  assign nw00304 = nw04263 ? \nr00026 [24] : nw00218;
  assign nw00305 = nw04263 ? \nr00026 [25] : nw00219;
  assign nw00306 = nw04263 ? \nr00026 [26] : nw00220;
  assign nw00307 = nw04263 ? \nr00026 [27] : nw00221;
  assign nw00308 = nw04263 ? \nr00026 [28] : nw00222;
  assign nw00309 = nw04263 ? \nr00026 [29] : nw00223;
  assign nw00310 = nw04263 ? \nr00026 [30] : nw00225;
  assign nw00311 = nw04263 ? \nr00026 [31] : nw00226;
  assign nw04269 = nw01388 & nw00455;
  assign nw04270 = nw00460 ? nw01388 : nw04269;
  assign nw00138 = nw04270 & ~(nw00454);
  assign nw04271 = ~(nw01416 & nw00455);
  assign nw04272 = nw00460 ? nw03284 : nw04271;
  assign nw00149 = \nr00025 [4] & ~(nw04272);
  assign nw04273 = ~\nr00066 [2];
  assign nw04274 = nw01444 & nw00455;
  assign nw04275 = nw00460 ? nw01444 : nw04274;
  assign nw00160 = \nr00025 [4] ? nw04275 : nw04273;
  assign nw04276 = \nr00066 [3] ^ \nr00066 [2];
  assign nw04277 = nw01472 & nw00455;
  assign nw04278 = nw00460 ? nw01472 : nw04277;
  assign nw00163 = \nr00025 [4] ? nw04278 : nw04276;
  assign nw04279 = \nr00066 [3] & \nr00066 [2];
  assign nw04280 = nw04279 ^ \nr00066 [4];
  assign nw04281 = nw01500 & nw00455;
  assign nw04282 = nw00460 ? nw01500 : nw04281;
  assign nw00164 = \nr00025 [4] ? nw04282 : nw04280;
  assign nw04283 = nw04279 & \nr00066 [4];
  assign nw04284 = nw04283 ^ \nr00066 [5];
  assign nw04285 = nw01528 & nw00455;
  assign nw04286 = nw00460 ? nw01528 : nw04285;
  assign nw00165 = \nr00025 [4] ? nw04286 : nw04284;
  assign nw04287 = ~(\nr00066 [5] & \nr00066 [4]);
  assign nw04288 = nw04279 & ~(nw04287);
  assign nw04289 = nw04288 ^ \nr00066 [6];
  assign nw04290 = nw01556 & nw00455;
  assign nw04291 = nw00460 ? nw01556 : nw04290;
  assign nw00166 = \nr00025 [4] ? nw04291 : nw04289;
  assign nw04292 = nw04288 & \nr00066 [6];
  assign nw04293 = nw04292 ^ \nr00066 [7];
  assign nw04294 = nw01584 & nw00455;
  assign nw04295 = nw00460 ? nw01584 : nw04294;
  assign nw00167 = \nr00025 [4] ? nw04295 : nw04293;
  assign nw04296 = ~(\nr00066 [7] & \nr00066 [6]);
  assign nw04297 = nw04288 & ~(nw04296);
  assign nw04298 = nw04297 ^ \nr00066 [8];
  assign nw04299 = nw01620 & nw00455;
  assign nw04300 = nw00460 ? nw01620 : nw04299;
  assign nw00168 = \nr00025 [4] ? nw04300 : nw04298;
  assign nw04301 = nw04297 & ~(nw01593);
  assign nw04302 = nw04301 ^ \nr00066 [9];
  assign nw04303 = nw01653 & nw00455;
  assign nw04304 = nw00460 ? nw01653 : nw04303;
  assign nw00169 = \nr00025 [4] ? nw04304 : nw04302;
  assign nw04305 = ~(\nr00066 [9] & \nr00066 [8]);
  assign nw04306 = nw04305 | nw04296;
  assign nw04307 = nw04288 & ~(nw04306);
  assign nw04308 = nw04307 ^ \nr00066 [10];
  assign nw04309 = nw01686 & nw00455;
  assign nw04310 = nw00460 ? nw01686 : nw04309;
  assign nw00139 = \nr00025 [4] ? nw04310 : nw04308;
  assign nw04311 = nw04307 & ~(nw01659);
  assign nw04312 = nw04311 ^ \nr00066 [11];
  assign nw04313 = nw01719 & nw00455;
  assign nw04314 = nw00460 ? nw01719 : nw04313;
  assign nw00140 = \nr00025 [4] ? nw04314 : nw04312;
  assign nw04315 = ~(\nr00066 [11] & \nr00066 [10]);
  assign nw04316 = nw04307 & ~(nw04315);
  assign nw04317 = nw04316 ^ \nr00066 [12];
  assign nw04318 = nw01752 & nw00455;
  assign nw04319 = nw00460 ? nw01752 : nw04318;
  assign nw00141 = \nr00025 [4] ? nw04319 : nw04317;
  assign nw04320 = nw04316 & ~(nw01725);
  assign nw04321 = nw04320 ^ \nr00066 [13];
  assign nw04322 = nw01785 & nw00455;
  assign nw04323 = nw00460 ? nw01785 : nw04322;
  assign nw00142 = \nr00025 [4] ? nw04323 : nw04321;
  assign nw04324 = ~(\nr00066 [13] & \nr00066 [12]);
  assign nw04325 = nw04324 | nw04315;
  assign nw04326 = nw04307 & ~(nw04325);
  assign nw04327 = nw04326 ^ \nr00066 [14];
  assign nw04328 = nw01818 & nw00455;
  assign nw04329 = nw00460 ? nw01818 : nw04328;
  assign nw00143 = \nr00025 [4] ? nw04329 : nw04327;
  assign nw04330 = nw04326 & ~(nw01791);
  assign nw04331 = nw04330 ^ \nr00066 [15];
  assign nw04332 = nw01849 & nw00455;
  assign nw04333 = nw00460 ? nw01849 : nw04332;
  assign nw00144 = \nr00025 [4] ? nw04333 : nw04331;
  assign nw04334 = ~(\nr00066 [15] & \nr00066 [14]);
  assign nw04335 = nw04326 & ~(nw04334);
  assign nw04336 = nw04335 ^ \nr00066 [16];
  assign nw04337 = nw01879 & nw00455;
  assign nw04338 = nw00460 ? nw01879 : nw04337;
  assign nw00145 = \nr00025 [4] ? nw04338 : nw04336;
  assign nw04339 = nw04335 & ~(nw01852);
  assign nw04340 = nw04339 ^ \nr00066 [17];
  assign nw04341 = nw01909 & nw00455;
  assign nw04342 = nw00460 ? nw01909 : nw04341;
  assign nw00146 = \nr00025 [4] ? nw04342 : nw04340;
  assign nw04343 = ~(\nr00066 [17] & \nr00066 [16]);
  assign nw04344 = nw04343 | nw04334;
  assign nw04345 = nw04344 | nw04325;
  assign nw04346 = nw04307 & ~(nw04345);
  assign nw04347 = nw04346 ^ \nr00066 [18];
  assign nw04348 = nw01939 & nw00455;
  assign nw04349 = nw00460 ? nw01939 : nw04348;
  assign nw00147 = \nr00025 [4] ? nw04349 : nw04347;
  assign nw04350 = nw04346 & ~(nw01912);
  assign nw04351 = nw04350 ^ \nr00066 [19];
  assign nw04352 = nw01969 & nw00455;
  assign nw04353 = nw00460 ? nw01969 : nw04352;
  assign nw00148 = \nr00025 [4] ? nw04353 : nw04351;
  assign nw04354 = ~(\nr00066 [19] & \nr00066 [18]);
  assign nw04355 = nw04346 & ~(nw04354);
  assign nw04356 = nw04355 ^ \nr00066 [20];
  assign nw04357 = nw01999 & nw00455;
  assign nw04358 = nw00460 ? nw01999 : nw04357;
  assign nw00150 = \nr00025 [4] ? nw04358 : nw04356;
  assign nw04359 = nw04355 & ~(nw01972);
  assign nw04360 = nw04359 ^ \nr00066 [21];
  assign nw04361 = nw02029 & nw00455;
  assign nw04362 = nw00460 ? nw02029 : nw04361;
  assign nw00151 = \nr00025 [4] ? nw04362 : nw04360;
  assign nw04363 = ~(\nr00066 [21] & \nr00066 [20]);
  assign nw04364 = nw04363 | nw04354;
  assign nw04365 = nw04346 & ~(nw04364);
  assign nw04366 = nw04365 ^ \nr00066 [22];
  assign nw04367 = nw02059 & nw00455;
  assign nw04368 = nw00460 ? nw02059 : nw04367;
  assign nw00152 = \nr00025 [4] ? nw04368 : nw04366;
  assign nw04369 = nw04365 & ~(nw02032);
  assign nw04370 = nw04369 ^ \nr00066 [23];
  assign nw04371 = nw02088 & nw00455;
  assign nw04372 = nw00460 ? nw02088 : nw04371;
  assign nw00153 = \nr00025 [4] ? nw04372 : nw04370;
  assign nw04373 = ~(\nr00066 [23] & \nr00066 [22]);
  assign nw04374 = nw04365 & ~(nw04373);
  assign nw04375 = nw04374 ^ \nr00066 [24];
  assign nw04376 = nw02117 & nw00455;
  assign nw04377 = nw00460 ? nw02117 : nw04376;
  assign nw00154 = \nr00025 [4] ? nw04377 : nw04375;
  assign nw04378 = nw04374 & ~(nw02090);
  assign nw04379 = nw04378 ^ \nr00066 [25];
  assign nw04380 = nw02146 & nw00455;
  assign nw04381 = nw00460 ? nw02146 : nw04380;
  assign nw00155 = \nr00025 [4] ? nw04381 : nw04379;
  assign nw04382 = ~(\nr00066 [25] & \nr00066 [24]);
  assign nw04383 = nw04382 | nw04373;
  assign nw04384 = nw04383 | nw04364;
  assign nw04385 = nw04346 & ~(nw04384);
  assign nw04386 = nw04385 ^ \nr00066 [26];
  assign nw04387 = nw02175 & nw00455;
  assign nw04388 = nw00460 ? nw02175 : nw04387;
  assign nw00156 = \nr00025 [4] ? nw04388 : nw04386;
  assign nw04389 = nw04385 & ~(nw02148);
  assign nw04390 = nw04389 ^ \nr00066 [27];
  assign nw04391 = nw02204 & nw00455;
  assign nw04392 = nw00460 ? nw02204 : nw04391;
  assign nw00157 = \nr00025 [4] ? nw04392 : nw04390;
  assign nw04393 = ~(\nr00066 [27] & \nr00066 [26]);
  assign nw04394 = nw04385 & ~(nw04393);
  assign nw04395 = nw04394 ^ \nr00066 [28];
  assign nw04396 = nw02233 & nw00455;
  assign nw04397 = nw00460 ? nw02233 : nw04396;
  assign nw00158 = \nr00025 [4] ? nw04397 : nw04395;
  assign nw04398 = nw04394 & ~(nw02206);
  assign nw04399 = nw04398 ^ \nr00066 [29];
  assign nw04400 = nw02262 & nw00455;
  assign nw04401 = nw00460 ? nw02262 : nw04400;
  assign nw00159 = \nr00025 [4] ? nw04401 : nw04399;
  assign nw04402 = ~(\nr00066 [29] & \nr00066 [28]);
  assign nw04403 = nw04402 | nw04393;
  assign nw04404 = nw04385 & ~(nw04403);
  assign nw04405 = nw04404 ^ \nr00066 [30];
  assign nw04406 = nw02291 & nw00455;
  assign nw04407 = nw00460 ? nw02291 : nw04406;
  assign nw00161 = \nr00025 [4] ? nw04407 : nw04405;
  assign nw04408 = nw04404 & ~(nw02264);
  assign nw04409 = nw04408 ^ \nr00066 [31];
  assign nw04410 = nw02320 & nw00455;
  assign nw04411 = nw00460 ? nw02320 : nw04410;
  assign nw00162 = \nr00025 [4] ? nw04411 : nw04409;
  assign nw04412 = nw01416 & ~(nw01388);
  assign nw04413 = nw04412 ? nw00202 : nw00209;
  assign nw04414 = \nr00048  ? nw04413 : nw00209;
  assign nw04415 = nw01416 ? nw00202 : nw04414;
  assign nw04416 = \nr00049  ? nw04415 : nw04414;
  assign nw00282 = \nr00060  ? nw00209 : nw04416;
  assign nw04417 = nw04412 ? nw00213 : nw00210;
  assign nw04418 = \nr00048  ? nw04417 : nw00210;
  assign nw04419 = nw01416 ? nw00213 : nw04418;
  assign nw04420 = \nr00049  ? nw04419 : nw04418;
  assign nw00283 = \nr00060  ? nw00210 : nw04420;
  assign nw04421 = nw04412 ? nw00224 : nw00211;
  assign nw04422 = \nr00048  ? nw04421 : nw00211;
  assign nw04423 = nw01416 ? nw00224 : nw04422;
  assign nw04424 = \nr00049  ? nw04423 : nw04422;
  assign nw00284 = \nr00060  ? nw00211 : nw04424;
  assign nw04425 = nw04412 ? nw00227 : nw00212;
  assign nw04426 = \nr00048  ? nw04425 : nw00212;
  assign nw04427 = nw01416 ? nw00227 : nw04426;
  assign nw04428 = \nr00049  ? nw04427 : nw04426;
  assign nw00285 = \nr00060  ? nw00212 : nw04428;
  assign nw04429 = nw04412 ? nw00228 : nw00214;
  assign nw04430 = \nr00048  ? nw04429 : nw00214;
  assign nw04431 = nw01416 ? nw00228 : nw04430;
  assign nw04432 = \nr00049  ? nw04431 : nw04430;
  assign nw00286 = \nr00060  ? nw00214 : nw04432;
  assign nw04433 = nw04412 ? nw00229 : nw00215;
  assign nw04434 = \nr00048  ? nw04433 : nw00215;
  assign nw04435 = nw01416 ? nw00229 : nw04434;
  assign nw04436 = \nr00049  ? nw04435 : nw04434;
  assign nw00287 = \nr00060  ? nw00215 : nw04436;
  assign nw04437 = nw04412 ? nw00230 : nw00216;
  assign nw04438 = \nr00048  ? nw04437 : nw00216;
  assign nw04439 = nw01416 ? nw00230 : nw04438;
  assign nw04440 = \nr00049  ? nw04439 : nw04438;
  assign nw00288 = \nr00060  ? nw00216 : nw04440;
  assign nw04441 = nw04412 ? nw00231 : nw00217;
  assign nw04442 = \nr00048  ? nw04441 : nw00217;
  assign nw04443 = nw01416 ? nw00231 : nw04442;
  assign nw04444 = \nr00049  ? nw04443 : nw04442;
  assign nw00289 = \nr00060  ? nw00217 : nw04444;
  assign nw04445 = nw01388 & ~(nw01416);
  assign nw04446 = nw04445 ? nw00202 : nw00232;
  assign nw04447 = \nr00048  ? nw04446 : nw00232;
  assign nw04448 = nw01416 ? nw04447 : nw00232;
  assign nw04449 = \nr00049  ? nw04448 : nw04447;
  assign nw00274 = \nr00060  ? nw00232 : nw04449;
  assign nw04450 = nw04445 ? nw00213 : nw00233;
  assign nw04451 = \nr00048  ? nw04450 : nw00233;
  assign nw04452 = nw01416 ? nw04451 : nw00233;
  assign nw04453 = \nr00049  ? nw04452 : nw04451;
  assign nw00275 = \nr00060  ? nw00233 : nw04453;
  assign nw04454 = nw04445 ? nw00224 : nw00203;
  assign nw04455 = \nr00048  ? nw04454 : nw00203;
  assign nw04456 = nw01416 ? nw04455 : nw00203;
  assign nw04457 = \nr00049  ? nw04456 : nw04455;
  assign nw00276 = \nr00060  ? nw00203 : nw04457;
  assign nw04458 = nw04445 ? nw00227 : nw00204;
  assign nw04459 = \nr00048  ? nw04458 : nw00204;
  assign nw04460 = nw01416 ? nw04459 : nw00204;
  assign nw04461 = \nr00049  ? nw04460 : nw04459;
  assign nw00277 = \nr00060  ? nw00204 : nw04461;
  assign nw04462 = nw04445 ? nw00228 : nw00205;
  assign nw04463 = \nr00048  ? nw04462 : nw00205;
  assign nw04464 = nw01416 ? nw04463 : nw00205;
  assign nw04465 = \nr00049  ? nw04464 : nw04463;
  assign nw00278 = \nr00060  ? nw00205 : nw04465;
  assign nw04466 = nw04445 ? nw00229 : nw00206;
  assign nw04467 = \nr00048  ? nw04466 : nw00206;
  assign nw04468 = nw01416 ? nw04467 : nw00206;
  assign nw04469 = \nr00049  ? nw04468 : nw04467;
  assign nw00279 = \nr00060  ? nw00206 : nw04469;
  assign nw04470 = nw04445 ? nw00230 : nw00207;
  assign nw04471 = \nr00048  ? nw04470 : nw00207;
  assign nw04472 = nw01416 ? nw04471 : nw00207;
  assign nw04473 = \nr00049  ? nw04472 : nw04471;
  assign nw00280 = \nr00060  ? nw00207 : nw04473;
  assign nw04474 = nw04445 ? nw00231 : nw00208;
  assign nw04475 = \nr00048  ? nw04474 : nw00208;
  assign nw04476 = nw01416 ? nw04475 : nw00208;
  assign nw04477 = \nr00049  ? nw04476 : nw04475;
  assign nw00281 = \nr00060  ? nw00208 : nw04477;
  assign nw04478 = nw01416 & nw01388;
  assign nw04479 = nw04478 ? nw00202 : nw00218;
  assign nw04480 = \nr00048  ? nw04479 : nw00218;
  assign nw04481 = nw01416 ? nw00232 : nw04480;
  assign nw04482 = \nr00049  ? nw04481 : nw04480;
  assign nw00266 = \nr00060  ? nw00218 : nw04482;
  assign nw04483 = nw04478 ? nw00213 : nw00219;
  assign nw04484 = \nr00048  ? nw04483 : nw00219;
  assign nw04485 = nw01416 ? nw00233 : nw04484;
  assign nw04486 = \nr00049  ? nw04485 : nw04484;
  assign nw00267 = \nr00060  ? nw00219 : nw04486;
  assign nw04487 = nw04478 ? nw00224 : nw00220;
  assign nw04488 = \nr00048  ? nw04487 : nw00220;
  assign nw04489 = nw01416 ? nw00203 : nw04488;
  assign nw04490 = \nr00049  ? nw04489 : nw04488;
  assign nw00268 = \nr00060  ? nw00220 : nw04490;
  assign nw04491 = nw04478 ? nw00227 : nw00221;
  assign nw04492 = \nr00048  ? nw04491 : nw00221;
  assign nw04493 = nw01416 ? nw00204 : nw04492;
  assign nw04494 = \nr00049  ? nw04493 : nw04492;
  assign nw00269 = \nr00060  ? nw00221 : nw04494;
  assign nw04495 = nw04478 ? nw00228 : nw00222;
  assign nw04496 = \nr00048  ? nw04495 : nw00222;
  assign nw04497 = nw01416 ? nw00205 : nw04496;
  assign nw04498 = \nr00049  ? nw04497 : nw04496;
  assign nw00270 = \nr00060  ? nw00222 : nw04498;
  assign nw04499 = nw04478 ? nw00229 : nw00223;
  assign nw04500 = \nr00048  ? nw04499 : nw00223;
  assign nw04501 = nw01416 ? nw00206 : nw04500;
  assign nw04502 = \nr00049  ? nw04501 : nw04500;
  assign nw00271 = \nr00060  ? nw00223 : nw04502;
  assign nw04503 = nw04478 ? nw00230 : nw00225;
  assign nw04504 = \nr00048  ? nw04503 : nw00225;
  assign nw04505 = nw01416 ? nw00207 : nw04504;
  assign nw04506 = \nr00049  ? nw04505 : nw04504;
  assign nw00272 = \nr00060  ? nw00225 : nw04506;
  assign nw04507 = nw04478 ? nw00231 : nw00226;
  assign nw04508 = \nr00048  ? nw04507 : nw00226;
  assign nw04509 = nw01416 ? nw00208 : nw04508;
  assign nw04510 = \nr00049  ? nw04509 : nw04508;
  assign nw00273 = \nr00060  ? nw00226 : nw04510;
  assign nw04511 = ~\nr00103 [2];
  assign nw04512 = \nr00103 [0] & ~(\nr00103 [1]);
  assign nw04513 = ~(\nr00103 [1] | \nr00103 [0]);
  assign nw04514 = \nr00103 [2] ? nw04513 : nw04512;
  assign nw04515 = \nr00103 [1] & \nr00103 [0];
  assign nw04516 = \nr00103 [2] ? nw04512 : nw04515;
  assign segmentos_o[0] = \nr00103 [3] ? nw04516 : nw04514;
  assign nw04517 = \nr00103 [1] & ~(\nr00103 [0]);
  assign nw04518 = ~(nw04517 | nw04512);
  assign nw04519 = \nr00103 [2] & ~(nw04518);
  assign nw04520 = \nr00103 [0] ? \nr00103 [1] : \nr00103 [2];
  assign segmentos_o[1] = \nr00103 [3] ? nw04520 : nw04519;
  assign nw04521 = \nr00103 [2] & ~(nw04512);
  assign nw04522 = nw04517 & ~(\nr00103 [2]);
  assign segmentos_o[2] = \nr00103 [3] ? nw04521 : nw04522;
  assign nw04523 = nw04515 | nw04513;
  assign nw04524 = \nr00103 [2] ? nw04523 : nw04512;
  assign nw04525 = \nr00103 [2] ? nw04515 : nw04517;
  assign segmentos_o[3] = \nr00103 [3] ? nw04525 : nw04524;
  assign nw04526 = nw04512 & ~(\nr00103 [2]);
  assign nw04527 = \nr00103 [0] | ~(\nr00103 [1]);
  assign nw04528 = \nr00103 [2] ? nw04527 : \nr00103 [0];
  assign segmentos_o[4] = \nr00103 [3] ? nw04526 : nw04528;
  assign nw04529 = nw04512 & ~(nw04511);
  assign nw04530 = \nr00103 [1] | \nr00103 [0];
  assign nw04531 = \nr00103 [2] ? nw04515 : nw04530;
  assign segmentos_o[5] = \nr00103 [3] ? nw04529 : nw04531;
  assign nw04532 = nw04513 & ~(nw04511);
  assign nw04533 = ~\nr00103 [1];
  assign nw04534 = \nr00103 [2] ? nw04515 : nw04533;
  assign segmentos_o[6] = \nr00103 [3] ? nw04532 : nw04534;
  assign nw04535 = ~\nw05427 [16];
  assign nw04536 = \nw05427 [15] | ~(\nw05427 [14]);
  assign nw04537 = nw04535 & ~(nw04536);
  assign nw04538 = nw04537 ? \nr00104 [4] : \nr00104 [0];
  assign nw04539 = ~(\nw05427 [15] & \nw05427 [14]);
  assign nw04540 = nw04539 | nw04535;
  assign nw04541 = \nw05427 [14] | ~(\nw05427 [15]);
  assign nw04542 = \nw05427 [16] & ~(nw04541);
  assign nw04543 = nw04540 & ~(nw04542);
  assign nw04544 = \nw05427 [16] & ~(nw04536);
  assign nw04545 = \nw05427 [15] | \nw05427 [14];
  assign nw04546 = \nw05427 [16] & ~(nw04545);
  assign nw04547 = nw04546 | nw04544;
  assign nw04548 = nw04543 & ~(nw04547);
  assign nw04549 = nw04535 & ~(nw04539);
  assign nw04550 = nw04535 & ~(nw04541);
  assign nw04551 = nw04550 | nw04549;
  assign nw04552 = nw04548 & ~(nw04551);
  assign nw04553 = \nr00104 [28] & ~(nw04540);
  assign nw04554 = nw04542 & \nr00104 [24];
  assign nw04555 = nw04554 | nw04553;
  assign nw04556 = nw04544 & \nr00104 [20];
  assign nw04557 = nw04546 & \nr00104 [16];
  assign nw04558 = nw04557 | nw04556;
  assign nw04559 = nw04558 | nw04555;
  assign nw04560 = nw04549 & \nr00104 [12];
  assign nw04561 = nw04550 & \nr00104 [8];
  assign nw04562 = nw04561 | nw04560;
  assign nw04563 = nw04562 | nw04559;
  assign nw05420[0] = nw04552 ? nw04538 : nw04563;
  assign nw04564 = nw04537 ? \nr00104 [5] : \nr00104 [1];
  assign nw04565 = nw04549 ? \nr00104 [13] : nw04564;
  assign nw04566 = ~(nw00882 & nw00418);
  assign nw04567 = nw04566 & ~(nw00434);
  assign nw04568 = nw00437 & ~(nw04567);
  assign nw04569 = ~(nw04568 | nw04565);
  assign nw04570 = ~nw04569;
  assign nw04571 = \nr00104 [29] & ~(nw04540);
  assign nw04572 = nw04542 & \nr00104 [25];
  assign nw04573 = nw04572 | nw04571;
  assign nw04574 = nw04544 & \nr00104 [21];
  assign nw04575 = nw04546 & \nr00104 [17];
  assign nw04576 = nw04575 | nw04574;
  assign nw04577 = nw04576 | nw04573;
  assign nw04578 = nw04549 & ~(nw04569);
  assign nw04579 = nw04550 & \nr00104 [9];
  assign nw04580 = nw04579 | nw04578;
  assign nw04581 = nw04580 | nw04577;
  assign nw05420[1] = nw04552 ? nw04570 : nw04581;
  assign nw04582 = nw04537 ? \nr00104 [6] : \nr00104 [2];
  assign nw04583 = \nr00104 [30] & ~(nw04540);
  assign nw04584 = nw04542 & \nr00104 [26];
  assign nw04585 = nw04584 | nw04583;
  assign nw04586 = nw04544 & \nr00104 [22];
  assign nw04587 = nw04546 & \nr00104 [18];
  assign nw04588 = nw04587 | nw04586;
  assign nw04589 = nw04588 | nw04585;
  assign nw04590 = nw04549 & \nr00104 [14];
  assign nw04591 = nw04550 & \nr00104 [10];
  assign nw04592 = nw04591 | nw04590;
  assign nw04593 = nw04592 | nw04589;
  assign nw05420[2] = nw04552 ? nw04582 : nw04593;
  assign nw04594 = nw04537 ? \nr00104 [7] : \nr00104 [3];
  assign nw04595 = \nr00104 [31] & ~(nw04540);
  assign nw04596 = nw04542 & \nr00104 [27];
  assign nw04597 = nw04596 | nw04595;
  assign nw04598 = nw04544 & \nr00104 [23];
  assign nw04599 = nw04546 & \nr00104 [19];
  assign nw04600 = nw04599 | nw04598;
  assign nw04601 = nw04600 | nw04597;
  assign nw04602 = nw04549 & \nr00104 [15];
  assign nw04603 = nw04550 & \nr00104 [11];
  assign nw04604 = nw04603 | nw04602;
  assign nw04605 = nw04604 | nw04601;
  assign nw05420[3] = nw04552 ? nw04594 : nw04605;
  assign nw04606 = ~(nw00102 | nw00103);
  assign nw04607 = nw04606 & ~(nw05416[0]);
  assign nw04608 = nw00957 | \nr00064 [6];
  assign nw04609 = nw04608 | nw00960;
  assign nw04610 = nw00960 | nw00958;
  assign nw04611 = ~(nw04610 & nw04609);
  assign nw04612 = nw04607 & ~(nw04611);
  assign nw04613 = \nr00064 [7] & ~(nw04609);
  assign nw05417[0] = nw04612 ? \nr00064 [20] : nw04613;
  assign nw04614 = nw05416[0] & ~(nw02000);
  assign nw04615 = \nr00064 [8] & ~(nw04610);
  assign nw04616 = \nr00064 [8] & ~(nw04609);
  assign nw04617 = nw04616 | nw04615;
  assign nw04618 = nw04617 | nw04614;
  assign nw05417[1] = nw04612 ? \nr00064 [21] : nw04618;
  assign nw04619 = nw05416[0] & ~(nw02030);
  assign nw04620 = \nr00064 [9] & ~(nw04610);
  assign nw04621 = \nr00064 [9] & ~(nw04609);
  assign nw04622 = nw04621 | nw04620;
  assign nw04623 = nw04622 | nw04619;
  assign nw05417[2] = nw04612 ? \nr00064 [22] : nw04623;
  assign nw04624 = nw05416[0] & ~(nw01590);
  assign nw04625 = \nr00064 [10] & ~(nw04610);
  assign nw04626 = \nr00064 [10] & ~(nw04609);
  assign nw04627 = nw04626 | nw04625;
  assign nw04628 = nw04627 | nw04624;
  assign nw05417[3] = nw04612 ? \nr00064 [23] : nw04628;
  assign nw04629 = nw05416[0] & ~(nw01586);
  assign nw04630 = \nr00064 [11] & ~(nw04610);
  assign nw04631 = \nr00064 [11] & ~(nw04609);
  assign nw04632 = nw04631 | nw04630;
  assign nw04633 = nw04632 | nw04629;
  assign nw05417[4] = nw04612 ? \nr00064 [24] : nw04633;
  assign nw04634 = nw05416[0] & ~(nw01621);
  assign nw04635 = \nr00064 [25] & ~(nw04610);
  assign nw04636 = \nr00064 [25] & ~(nw04609);
  assign nw04637 = nw04636 | nw04635;
  assign nw04638 = nw04637 | nw04634;
  assign nw05417[5] = nw04612 ? \nr00064 [25] : nw04638;
  assign nw04639 = nw05416[0] & ~(nw01654);
  assign nw04640 = \nr00064 [26] & ~(nw04610);
  assign nw04641 = \nr00064 [26] & ~(nw04609);
  assign nw04642 = nw04641 | nw04640;
  assign nw04643 = nw04642 | nw04639;
  assign nw05417[6] = nw04612 ? \nr00064 [26] : nw04643;
  assign nw04644 = nw05416[0] & ~(nw01687);
  assign nw04645 = \nr00064 [27] & ~(nw04610);
  assign nw04646 = \nr00064 [27] & ~(nw04609);
  assign nw04647 = nw04646 | nw04645;
  assign nw04648 = nw04647 | nw04644;
  assign nw05417[7] = nw04612 ? \nr00064 [27] : nw04648;
  assign nw04649 = nw05416[0] & ~(nw01721);
  assign nw04650 = \nr00064 [28] & ~(nw04610);
  assign nw04651 = \nr00064 [28] & ~(nw04609);
  assign nw04652 = nw04651 | nw04650;
  assign nw04653 = nw04652 | nw04649;
  assign nw05417[8] = nw04612 ? \nr00064 [28] : nw04653;
  assign nw04654 = nw05416[0] & ~(nw01754);
  assign nw04655 = \nr00064 [29] & ~(nw04610);
  assign nw04656 = \nr00064 [29] & ~(nw04609);
  assign nw04657 = nw04656 | nw04655;
  assign nw04658 = nw04657 | nw04654;
  assign nw05417[9] = nw04612 ? \nr00064 [29] : nw04658;
  assign nw04659 = nw05416[0] & ~(nw01787);
  assign nw04660 = \nr00064 [30] & ~(nw04610);
  assign nw04661 = \nr00064 [30] & ~(nw04609);
  assign nw04662 = nw04661 | nw04660;
  assign nw04663 = nw04662 | nw04659;
  assign nw05417[10] = nw04612 ? \nr00064 [30] : nw04663;
  assign nw04664 = nw05416[0] & ~(nw00978);
  assign nw04665 = \nr00064 [7] & ~(nw04610);
  assign nw04666 = \nr00064 [31] & ~(nw04609);
  assign nw04667 = nw04666 | nw04665;
  assign nw04668 = nw04667 | nw04664;
  assign nw05417[11] = nw04612 ? \nr00064 [31] : nw04668;
  assign nw04669 = nw05416[0] & ~(nw01970);
  assign nw04670 = \nr00064 [12] & ~(nw04606);
  assign nw04671 = nw04670 | nw04669;
  assign nw04672 = \nr00064 [31] & ~(nw04610);
  assign nw04673 = nw04672 | nw04666;
  assign nw04674 = nw04673 | nw04671;
  assign nw05417[12] = nw04612 ? \nr00064 [31] : nw04674;
  assign nw04675 = nw05416[0] & ~(nw01720);
  assign nw04676 = \nr00064 [13] & ~(nw04606);
  assign nw04677 = nw04676 | nw04675;
  assign nw04678 = nw04677 | nw04673;
  assign nw05417[13] = nw04612 ? \nr00064 [31] : nw04678;
  assign nw04679 = nw05416[0] & ~(nw01753);
  assign nw04680 = \nr00064 [14] & ~(nw04606);
  assign nw04681 = nw04680 | nw04679;
  assign nw04682 = nw04681 | nw04673;
  assign nw05417[14] = nw04612 ? \nr00064 [31] : nw04682;
  assign nw04683 = nw05416[0] & ~(nw01786);
  assign nw04684 = \nr00064 [15] & ~(nw04606);
  assign nw04685 = nw04684 | nw04683;
  assign nw04686 = nw04685 | nw04673;
  assign nw05417[15] = nw04612 ? \nr00064 [31] : nw04686;
  assign nw04687 = nw05416[0] & ~(nw01591);
  assign nw04688 = \nr00064 [16] & ~(nw04606);
  assign nw04689 = nw04688 | nw04687;
  assign nw04690 = nw04689 | nw04673;
  assign nw05417[16] = nw04612 ? \nr00064 [31] : nw04690;
  assign nw04691 = nw05416[0] & ~(nw01850);
  assign nw04692 = \nr00064 [17] & ~(nw04606);
  assign nw04693 = nw04692 | nw04691;
  assign nw04694 = nw04693 | nw04673;
  assign nw05417[17] = nw04612 ? \nr00064 [31] : nw04694;
  assign nw04695 = nw05416[0] & ~(nw01880);
  assign nw04696 = \nr00064 [18] & ~(nw04606);
  assign nw04697 = nw04696 | nw04695;
  assign nw04698 = nw04697 | nw04673;
  assign nw05417[18] = nw04612 ? \nr00064 [31] : nw04698;
  assign nw04699 = nw05416[0] & ~(nw01910);
  assign nw04700 = \nr00064 [19] & ~(nw04606);
  assign nw04701 = nw04700 | nw04699;
  assign nw04702 = nw04701 | nw04673;
  assign nw05417[19] = nw04612 ? \nr00064 [31] : nw04702;
  assign nw04703 = nw05416[0] & ~(nw01940);
  assign nw04704 = \nr00064 [20] & ~(nw04606);
  assign nw04705 = nw04704 | nw04703;
  assign nw04706 = nw04705 | nw04673;
  assign nw05417[20] = nw04612 ? \nr00064 [31] : nw04706;
  assign nw04707 = \nr00064 [21] & ~(nw04606);
  assign nw04708 = nw04707 | nw04664;
  assign nw04709 = nw04708 | nw04673;
  assign nw05417[21] = nw04612 ? \nr00064 [31] : nw04709;
  assign nw04710 = \nr00064 [22] & ~(nw04606);
  assign nw04711 = nw04710 | nw04664;
  assign nw04712 = nw04711 | nw04673;
  assign nw05417[22] = nw04612 ? \nr00064 [31] : nw04712;
  assign nw04713 = \nr00064 [23] & ~(nw04606);
  assign nw04714 = nw04713 | nw04664;
  assign nw04715 = nw04714 | nw04673;
  assign nw05417[23] = nw04612 ? \nr00064 [31] : nw04715;
  assign nw04716 = \nr00064 [24] & ~(nw04606);
  assign nw04717 = nw04716 | nw04664;
  assign nw04718 = nw04717 | nw04673;
  assign nw05417[24] = nw04612 ? \nr00064 [31] : nw04718;
  assign nw04719 = \nr00064 [25] & ~(nw04606);
  assign nw04720 = nw04719 | nw04664;
  assign nw04721 = nw04720 | nw04673;
  assign nw05417[25] = nw04612 ? \nr00064 [31] : nw04721;
  assign nw04722 = \nr00064 [26] & ~(nw04606);
  assign nw04723 = nw04722 | nw04664;
  assign nw04724 = nw04723 | nw04673;
  assign nw05417[26] = nw04612 ? \nr00064 [31] : nw04724;
  assign nw04725 = \nr00064 [27] & ~(nw04606);
  assign nw04726 = nw04725 | nw04664;
  assign nw04727 = nw04726 | nw04673;
  assign nw05417[27] = nw04612 ? \nr00064 [31] : nw04727;
  assign nw04728 = \nr00064 [28] & ~(nw04606);
  assign nw04729 = nw04728 | nw04664;
  assign nw04730 = nw04729 | nw04673;
  assign nw05417[28] = nw04612 ? \nr00064 [31] : nw04730;
  assign nw04731 = \nr00064 [29] & ~(nw04606);
  assign nw04732 = nw04731 | nw04664;
  assign nw04733 = nw04732 | nw04673;
  assign nw05417[29] = nw04612 ? \nr00064 [31] : nw04733;
  assign nw04734 = \nr00064 [30] & ~(nw04606);
  assign nw04735 = nw04734 | nw04664;
  assign nw04736 = nw04735 | nw04673;
  assign nw05417[30] = nw04612 ? \nr00064 [31] : nw04736;
  assign nw04737 = nw04535 & ~(nw04545);
  assign nw04738 = ~\nw05427 [14];
  assign nw04739 = ~(nw04737 & nw04738);
  assign nw04740 = nw04541 & nw04536;
  assign nw04741 = ~nw04740;
  assign nw04742 = nw04741 | nw04739;
  assign nw04743 = nw04545 ^ nw04535;
  assign nw04744 = nw04743 & ~(nw04742);
  assign anodos_o[0] = ~(nw04744 & nw04737);
  assign nw04745 = nw04737 | nw04738;
  assign nw04746 = nw04745 | nw04740;
  assign nw04747 = nw04746 | nw04743;
  assign anodos_o[1] = nw04747 | nw04737;
  assign nw04748 = nw04737 | \nw05427 [14];
  assign nw04749 = nw04748 | nw04740;
  assign nw04750 = nw04749 | nw04743;
  assign anodos_o[2] = nw04750 | nw04737;
  assign nw04751 = nw04745 | nw04741;
  assign nw04752 = nw04751 | nw04743;
  assign anodos_o[3] = nw04752 | nw04737;
  assign nw04753 = nw04748 | nw04741;
  assign nw04754 = nw04753 | nw04743;
  assign anodos_o[4] = nw04754 | nw04737;
  assign nw04755 = ~nw04743;
  assign nw04756 = nw04746 | nw04755;
  assign anodos_o[5] = nw04756 | nw04737;
  assign nw04757 = nw04749 | nw04755;
  assign anodos_o[6] = nw04757 | nw04737;
  assign nw04758 = nw04751 | nw04755;
  assign anodos_o[7] = nw04758 | nw04737;
  assign nw04759 = \nr00016 [31] & ~(\nr00017 [31]);
  assign nw00258 = \nr00016 [31] | \nr00017 [31];
  assign nw05413[31] = \nr00016 [31] & \nr00017 [31];
  assign nw04760 = nw00258 & ~(nw05413[31]);
  assign nw04761 = \nr00017 [30] | ~(\nr00016 [30]);
  assign nw04762 = ~(nw04761 | nw04760);
  assign nw04763 = ~(nw04762 | nw04759);
  assign nw00257 = \nr00016 [30] | \nr00017 [30];
  assign nw05413[30] = \nr00016 [30] & \nr00017 [30];
  assign nw04764 = nw00257 & ~(nw05413[30]);
  assign nw04765 = ~(nw04764 | nw04760);
  assign nw04766 = \nr00017 [29] | ~(\nr00016 [29]);
  assign nw00255 = \nr00016 [29] | \nr00017 [29];
  assign nw05413[29] = \nr00016 [29] & \nr00017 [29];
  assign nw04767 = nw00255 & ~(nw05413[29]);
  assign nw04768 = \nr00017 [28] | ~(\nr00016 [28]);
  assign nw04769 = ~(nw04768 | nw04767);
  assign nw04770 = nw04766 & ~(nw04769);
  assign nw04771 = nw04765 & ~(nw04770);
  assign nw04772 = nw04763 & ~(nw04771);
  assign nw00254 = \nr00016 [28] | \nr00017 [28];
  assign nw05413[28] = \nr00016 [28] & \nr00017 [28];
  assign nw04773 = nw00254 & ~(nw05413[28]);
  assign nw04774 = ~(nw04773 | nw04767);
  assign nw04775 = nw04774 & nw04765;
  assign nw04776 = \nr00017 [27] | ~(\nr00016 [27]);
  assign nw00253 = \nr00016 [27] | \nr00017 [27];
  assign nw05413[27] = \nr00016 [27] & \nr00017 [27];
  assign nw04777 = nw00253 & ~(nw05413[27]);
  assign nw04778 = \nr00017 [26] | ~(\nr00016 [26]);
  assign nw04779 = ~(nw04778 | nw04777);
  assign nw04780 = nw04776 & ~(nw04779);
  assign nw00252 = \nr00016 [26] | \nr00017 [26];
  assign nw05413[26] = \nr00016 [26] & \nr00017 [26];
  assign nw04781 = nw00252 & ~(nw05413[26]);
  assign nw04782 = ~(nw04781 | nw04777);
  assign nw04783 = \nr00017 [25] | ~(\nr00016 [25]);
  assign nw00251 = \nr00016 [25] | \nr00017 [25];
  assign nw05413[25] = \nr00016 [25] & \nr00017 [25];
  assign nw04784 = nw00251 & ~(nw05413[25]);
  assign nw04785 = \nr00017 [24] | ~(\nr00016 [24]);
  assign nw04786 = ~(nw04785 | nw04784);
  assign nw04787 = nw04783 & ~(nw04786);
  assign nw04788 = nw04782 & ~(nw04787);
  assign nw04789 = nw04780 & ~(nw04788);
  assign nw04790 = nw04775 & ~(nw04789);
  assign nw04791 = nw04772 & ~(nw04790);
  assign nw00250 = \nr00016 [24] | \nr00017 [24];
  assign nw05413[24] = \nr00016 [24] & \nr00017 [24];
  assign nw04792 = nw00250 & ~(nw05413[24]);
  assign nw04793 = ~(nw04792 | nw04784);
  assign nw04794 = nw04793 & nw04782;
  assign nw04795 = nw04794 & nw04775;
  assign nw04796 = \nr00017 [23] | ~(\nr00016 [23]);
  assign nw00249 = \nr00016 [23] | \nr00017 [23];
  assign nw05413[23] = \nr00016 [23] & \nr00017 [23];
  assign nw04797 = nw00249 & ~(nw05413[23]);
  assign nw04798 = \nr00017 [22] | ~(\nr00016 [22]);
  assign nw04799 = ~(nw04798 | nw04797);
  assign nw04800 = nw04796 & ~(nw04799);
  assign nw00248 = \nr00016 [22] | \nr00017 [22];
  assign nw05413[22] = \nr00016 [22] & \nr00017 [22];
  assign nw04801 = nw00248 & ~(nw05413[22]);
  assign nw04802 = ~(nw04801 | nw04797);
  assign nw04803 = \nr00017 [21] | ~(\nr00016 [21]);
  assign nw00247 = \nr00016 [21] | \nr00017 [21];
  assign nw05413[21] = \nr00016 [21] & \nr00017 [21];
  assign nw04804 = nw00247 & ~(nw05413[21]);
  assign nw04805 = \nr00017 [20] | ~(\nr00016 [20]);
  assign nw04806 = ~(nw04805 | nw04804);
  assign nw04807 = nw04803 & ~(nw04806);
  assign nw04808 = nw04802 & ~(nw04807);
  assign nw04809 = nw04800 & ~(nw04808);
  assign nw00246 = \nr00016 [20] | \nr00017 [20];
  assign nw05413[20] = \nr00016 [20] & \nr00017 [20];
  assign nw04810 = nw00246 & ~(nw05413[20]);
  assign nw04811 = ~(nw04810 | nw04804);
  assign nw04812 = nw04811 & nw04802;
  assign nw04813 = \nr00017 [19] | ~(\nr00016 [19]);
  assign nw00244 = \nr00016 [19] | \nr00017 [19];
  assign nw05413[19] = \nr00016 [19] & \nr00017 [19];
  assign nw04814 = nw00244 & ~(nw05413[19]);
  assign nw04815 = \nr00017 [18] | ~(\nr00016 [18]);
  assign nw04816 = ~(nw04815 | nw04814);
  assign nw04817 = nw04813 & ~(nw04816);
  assign nw00243 = \nr00016 [18] | \nr00017 [18];
  assign nw05413[18] = \nr00016 [18] & \nr00017 [18];
  assign nw04818 = nw00243 & ~(nw05413[18]);
  assign nw04819 = ~(nw04818 | nw04814);
  assign nw04820 = \nr00017 [17] | ~(\nr00016 [17]);
  assign nw00242 = \nr00016 [17] | \nr00017 [17];
  assign nw05413[17] = \nr00016 [17] & \nr00017 [17];
  assign nw04821 = nw00242 & ~(nw05413[17]);
  assign nw04822 = \nr00017 [16] | ~(\nr00016 [16]);
  assign nw04823 = ~(nw04822 | nw04821);
  assign nw04824 = nw04820 & ~(nw04823);
  assign nw04825 = nw04819 & ~(nw04824);
  assign nw04826 = nw04817 & ~(nw04825);
  assign nw04827 = nw04812 & ~(nw04826);
  assign nw04828 = nw04809 & ~(nw04827);
  assign nw04829 = nw04795 & ~(nw04828);
  assign nw04830 = nw04791 & ~(nw04829);
  assign nw00241 = \nr00016 [16] | \nr00017 [16];
  assign nw05413[16] = \nr00016 [16] & \nr00017 [16];
  assign nw04831 = nw00241 & ~(nw05413[16]);
  assign nw04832 = ~(nw04831 | nw04821);
  assign nw04833 = nw04832 & nw04819;
  assign nw04834 = nw04833 & nw04812;
  assign nw04835 = nw04834 & nw04795;
  assign nw04836 = \nr00017 [15] | ~(\nr00016 [15]);
  assign nw00240 = \nr00016 [15] | \nr00017 [15];
  assign nw05413[15] = \nr00016 [15] & \nr00017 [15];
  assign nw04837 = nw00240 & ~(nw05413[15]);
  assign nw04838 = \nr00017 [14] | ~(\nr00016 [14]);
  assign nw04839 = ~(nw04838 | nw04837);
  assign nw04840 = nw04836 & ~(nw04839);
  assign nw00239 = \nr00016 [14] | \nr00017 [14];
  assign nw05413[14] = \nr00016 [14] & \nr00017 [14];
  assign nw04841 = nw00239 & ~(nw05413[14]);
  assign nw04842 = ~(nw04841 | nw04837);
  assign nw04843 = \nr00017 [13] | ~(\nr00016 [13]);
  assign nw00238 = \nr00016 [13] | \nr00017 [13];
  assign nw05413[13] = \nr00016 [13] & \nr00017 [13];
  assign nw04844 = nw00238 & ~(nw05413[13]);
  assign nw04845 = \nr00017 [12] | ~(\nr00016 [12]);
  assign nw04846 = ~(nw04845 | nw04844);
  assign nw04847 = nw04843 & ~(nw04846);
  assign nw04848 = nw04842 & ~(nw04847);
  assign nw04849 = nw04840 & ~(nw04848);
  assign nw00237 = \nr00016 [12] | \nr00017 [12];
  assign nw05413[12] = \nr00016 [12] & \nr00017 [12];
  assign nw04850 = nw00237 & ~(nw05413[12]);
  assign nw04851 = ~(nw04850 | nw04844);
  assign nw04852 = nw04851 & nw04842;
  assign nw04853 = \nr00017 [11] | ~(\nr00016 [11]);
  assign nw00236 = \nr00016 [11] | \nr00017 [11];
  assign nw05413[11] = \nr00016 [11] & \nr00017 [11];
  assign nw04854 = nw00236 & ~(nw05413[11]);
  assign nw04855 = \nr00017 [10] | ~(\nr00016 [10]);
  assign nw04856 = ~(nw04855 | nw04854);
  assign nw04857 = nw04853 & ~(nw04856);
  assign nw00235 = \nr00016 [10] | \nr00017 [10];
  assign nw05413[10] = \nr00016 [10] & \nr00017 [10];
  assign nw04858 = nw00235 & ~(nw05413[10]);
  assign nw04859 = ~(nw04858 | nw04854);
  assign nw04860 = \nr00017 [9] | ~(\nr00016 [9]);
  assign nw00265 = \nr00016 [9] | \nr00017 [9];
  assign nw05413[9] = \nr00016 [9] & \nr00017 [9];
  assign nw04861 = nw00265 & ~(nw05413[9]);
  assign nw04862 = \nr00017 [8] | ~(\nr00016 [8]);
  assign nw04863 = ~(nw04862 | nw04861);
  assign nw04864 = nw04860 & ~(nw04863);
  assign nw04865 = nw04859 & ~(nw04864);
  assign nw04866 = nw04857 & ~(nw04865);
  assign nw04867 = nw04852 & ~(nw04866);
  assign nw04868 = nw04849 & ~(nw04867);
  assign nw00264 = \nr00016 [8] | \nr00017 [8];
  assign nw05413[8] = \nr00016 [8] & \nr00017 [8];
  assign nw04869 = nw00264 & ~(nw05413[8]);
  assign nw04870 = ~(nw04869 | nw04861);
  assign nw04871 = nw04870 & nw04859;
  assign nw04872 = nw04871 & nw04852;
  assign nw04873 = \nr00017 [7] | ~(\nr00016 [7]);
  assign nw00263 = \nr00016 [7] | \nr00017 [7];
  assign nw05413[7] = \nr00016 [7] & \nr00017 [7];
  assign nw04874 = nw00263 & ~(nw05413[7]);
  assign nw04875 = \nr00017 [6] | ~(\nr00016 [6]);
  assign nw04876 = ~(nw04875 | nw04874);
  assign nw04877 = nw04873 & ~(nw04876);
  assign nw00262 = \nr00016 [6] | \nr00017 [6];
  assign nw05413[6] = \nr00016 [6] & \nr00017 [6];
  assign nw04878 = nw00262 & ~(nw05413[6]);
  assign nw04879 = ~(nw04878 | nw04874);
  assign nw04880 = \nr00017 [5] | ~(\nr00016 [5]);
  assign nw00261 = \nr00016 [5] | \nr00017 [5];
  assign nw05413[5] = \nr00016 [5] & \nr00017 [5];
  assign nw04881 = nw00261 & ~(nw05413[5]);
  assign nw04882 = \nr00017 [4] | ~(\nr00016 [4]);
  assign nw04883 = ~(nw04882 | nw04881);
  assign nw04884 = nw04880 & ~(nw04883);
  assign nw04885 = nw04879 & ~(nw04884);
  assign nw04886 = nw04877 & ~(nw04885);
  assign nw00260 = \nr00016 [4] | \nr00017 [4];
  assign nw05413[4] = \nr00016 [4] & \nr00017 [4];
  assign nw04887 = nw00260 & ~(nw05413[4]);
  assign nw04888 = ~(nw04887 | nw04881);
  assign nw04889 = nw04888 & nw04879;
  assign nw04890 = \nr00017 [3] | ~(\nr00016 [3]);
  assign nw00259 = \nr00016 [3] | \nr00017 [3];
  assign nw05413[3] = \nr00016 [3] & \nr00017 [3];
  assign nw04891 = nw00259 & ~(nw05413[3]);
  assign nw04892 = \nr00017 [2] | ~(\nr00016 [2]);
  assign nw04893 = ~(nw04892 | nw04891);
  assign nw04894 = nw04890 & ~(nw04893);
  assign nw00256 = \nr00016 [2] | \nr00017 [2];
  assign nw05413[2] = \nr00016 [2] & \nr00017 [2];
  assign nw04895 = nw00256 & ~(nw05413[2]);
  assign nw04896 = ~(nw04895 | nw04891);
  assign nw04897 = \nr00017 [1] | ~(\nr00016 [1]);
  assign nw00245 = \nr00016 [1] | \nr00017 [1];
  assign nw05413[1] = \nr00016 [1] & \nr00017 [1];
  assign nw04898 = nw00245 & ~(nw05413[1]);
  assign nw04899 = \nr00017 [0] & ~(\nr00016 [0]);
  assign nw04900 = ~(nw04899 | nw04898);
  assign nw04901 = nw04897 & ~(nw04900);
  assign nw04902 = nw04896 & ~(nw04901);
  assign nw04903 = nw04894 & ~(nw04902);
  assign nw04904 = nw04889 & ~(nw04903);
  assign nw04905 = nw04886 & ~(nw04904);
  assign nw04906 = nw04872 & ~(nw04905);
  assign nw04907 = nw04868 & ~(nw04906);
  assign nw04908 = nw04835 & ~(nw04907);
  assign nw00050 = nw04830 & ~(nw04908);
  assign nw04909 = nw00882 & nw05430[1];
  assign nw04910 = nw00882 & nw05430[2];
  assign nw04911 = ~(nw04910 | nw04909);
  assign nw04912 = nw00437 & ~(nw04911);
  assign led_o[0] = nw04912 | \nr00105 [0];
  assign nw04913 = nw00436 & ~(nw04909);
  assign nw04914 = nw00437 & ~(nw04913);
  assign led_o[1] = nw04914 | \nr00105 [1];
  assign nw04915 = nw04910 & nw00437;
  assign led_o[2] = nw04915 | \nr00105 [2];
  assign led_o[3] = \nr00105 [3] | nw05430[0];
  assign led_o[4] = nw04915 | \nr00105 [4];
  assign led_o[5] = \nr00105 [5] | nw05430[0];
  assign led_o[6] = nw04912 | \nr00105 [6];
  assign led_o[7] = nw04914 | \nr00105 [7];
  assign led_o[8] = nw04912 | \nr00105 [8];
  assign led_o[9] = nw04914 | \nr00105 [9];
  assign led_o[10] = nw04915 | \nr00105 [10];
  assign led_o[11] = \nr00105 [11] | nw05430[0];
  assign led_o[12] = nw04915 | \nr00105 [12];
  assign led_o[13] = \nr00105 [13] | nw05430[0];
  assign led_o[14] = nw04912 | \nr00105 [14];
  assign led_o[15] = nw04914 | \nr00105 [15];
  assign ext_bus_we_o = nr00008 & ~(nw01176);
  assign ram_we_o = nw01199 & nr00008;
  assign nw04916 = nw04834 & ~(nw04907);
  assign nw04917 = nw04828 & ~(nw04916);
  assign nw04918 = nw04794 & ~(nw04917);
  assign nw04919 = nw04789 & ~(nw04918);
  assign nw04920 = nw04774 & ~(nw04919);
  assign nw04921 = nw04770 & ~(nw04920);
  assign nw04922 = ~(nw04921 | nw04764);
  assign nw04923 = nw04761 & ~(nw04922);
  assign nw04924 = ~(nw04923 ^ nw04760);
  assign nw05409[31] = ~nw04924;
  assign nw00054 = nw00050 ^ nw04760;
  assign nw04925 = nw00659 | nw00589;
  assign nw00384 = nw00594 & ~(nw04925);
  assign nw05409[1] = nw04899 ^ nw04898;
  assign nw05409[2] = nw04901 ^ nw04895;
  assign nw04926 = ~(nw04901 | nw04895);
  assign nw04927 = nw04892 & ~(nw04926);
  assign nw05409[3] = nw04927 ^ nw04891;
  assign nw05409[4] = nw04903 ^ nw04887;
  assign nw04928 = ~(nw04903 | nw04887);
  assign nw04929 = nw04882 & ~(nw04928);
  assign nw05409[5] = nw04929 ^ nw04881;
  assign nw04930 = nw04888 & ~(nw04903);
  assign nw04931 = nw04884 & ~(nw04930);
  assign nw05409[6] = nw04931 ^ nw04878;
  assign nw04932 = ~(nw04931 | nw04878);
  assign nw04933 = nw04875 & ~(nw04932);
  assign nw05409[7] = nw04933 ^ nw04874;
  assign nw05409[8] = nw04905 ^ nw04869;
  assign nw04934 = ~(nw04905 | nw04869);
  assign nw04935 = nw04862 & ~(nw04934);
  assign nw05409[9] = nw04935 ^ nw04861;
  assign nw04936 = nw04870 & ~(nw04905);
  assign nw04937 = nw04864 & ~(nw04936);
  assign nw05409[10] = nw04937 ^ nw04858;
  assign nw04938 = ~(nw04937 | nw04858);
  assign nw04939 = nw04855 & ~(nw04938);
  assign nw05409[11] = nw04939 ^ nw04854;
  assign nw04940 = nw04871 & ~(nw04905);
  assign nw04941 = nw04866 & ~(nw04940);
  assign nw05409[12] = nw04941 ^ nw04850;
  assign nw04942 = ~(nw04941 | nw04850);
  assign nw04943 = nw04845 & ~(nw04942);
  assign nw05409[13] = nw04943 ^ nw04844;
  assign nw04944 = nw04851 & ~(nw04941);
  assign nw04945 = nw04847 & ~(nw04944);
  assign nw05409[14] = nw04945 ^ nw04841;
  assign nw04946 = ~(nw04945 | nw04841);
  assign nw04947 = nw04838 & ~(nw04946);
  assign nw05409[15] = nw04947 ^ nw04837;
  assign nw05409[16] = nw04907 ^ nw04831;
  assign nw04948 = ~(nw04907 | nw04831);
  assign nw04949 = nw04822 & ~(nw04948);
  assign nw05409[17] = nw04949 ^ nw04821;
  assign nw04950 = nw04832 & ~(nw04907);
  assign nw04951 = nw04824 & ~(nw04950);
  assign nw05409[18] = nw04951 ^ nw04818;
  assign nw04952 = ~(nw04951 | nw04818);
  assign nw04953 = nw04815 & ~(nw04952);
  assign nw05409[19] = nw04953 ^ nw04814;
  assign nw04954 = nw04833 & ~(nw04907);
  assign nw04955 = nw04826 & ~(nw04954);
  assign nw05409[20] = nw04955 ^ nw04810;
  assign nw04956 = ~(nw04955 | nw04810);
  assign nw04957 = nw04805 & ~(nw04956);
  assign nw05409[21] = nw04957 ^ nw04804;
  assign nw04958 = nw04811 & ~(nw04955);
  assign nw04959 = nw04807 & ~(nw04958);
  assign nw05409[22] = nw04959 ^ nw04801;
  assign nw04960 = ~(nw04959 | nw04801);
  assign nw04961 = nw04798 & ~(nw04960);
  assign nw05409[23] = nw04961 ^ nw04797;
  assign nw05409[24] = nw04917 ^ nw04792;
  assign nw04962 = ~(nw04917 | nw04792);
  assign nw04963 = nw04785 & ~(nw04962);
  assign nw05409[25] = nw04963 ^ nw04784;
  assign nw04964 = nw04793 & ~(nw04917);
  assign nw04965 = nw04787 & ~(nw04964);
  assign nw05409[26] = nw04965 ^ nw04781;
  assign nw04966 = ~(nw04965 | nw04781);
  assign nw04967 = nw04778 & ~(nw04966);
  assign nw05409[27] = nw04967 ^ nw04777;
  assign nw05409[28] = nw04919 ^ nw04773;
  assign nw04968 = ~(nw04919 | nw04773);
  assign nw04969 = nw04768 & ~(nw04968);
  assign nw05409[29] = nw04969 ^ nw04767;
  assign nw05409[30] = nw04921 ^ nw04764;
  assign nw04970 = ~(\nr00016 [1] ^ \nr00017 [1]);
  assign nw05411[1] = ~nw04970;
  assign nw05412[1] = ~(nw04970 ^ nw05410[0]);
  assign nw04971 = ~(\nr00016 [2] ^ \nr00017 [2]);
  assign nw05411[2] = ~nw04971;
  assign nw04972 = nw05410[0] & ~(nw04970);
  assign nw04973 = ~(nw04972 | nw05413[1]);
  assign nw05412[2] = nw04973 ^ nw04971;
  assign nw04974 = ~(\nr00016 [3] ^ \nr00017 [3]);
  assign nw05411[3] = ~nw04974;
  assign nw04975 = nw04973 | nw04971;
  assign nw04976 = nw04975 & ~(nw05413[2]);
  assign nw05412[3] = nw04976 ^ nw04974;
  assign nw04977 = ~(\nr00016 [4] ^ \nr00017 [4]);
  assign nw05411[4] = ~nw04977;
  assign nw04978 = nw05413[2] & ~(nw04974);
  assign nw04979 = ~(nw04978 | nw05413[3]);
  assign nw04980 = ~(nw04974 | nw04971);
  assign nw04981 = nw04980 & ~(nw04973);
  assign nw04982 = nw04979 & ~(nw04981);
  assign nw05412[4] = nw04982 ^ nw04977;
  assign nw04983 = ~(\nr00016 [5] ^ \nr00017 [5]);
  assign nw05411[5] = ~nw04983;
  assign nw04984 = nw04982 | nw04977;
  assign nw04985 = nw04984 & ~(nw05413[4]);
  assign nw05412[5] = nw04985 ^ nw04983;
  assign nw04986 = ~(\nr00016 [6] ^ \nr00017 [6]);
  assign nw05411[6] = ~nw04986;
  assign nw04987 = nw05413[4] & ~(nw04983);
  assign nw04988 = ~(nw04987 | nw05413[5]);
  assign nw04989 = nw04983 | nw04977;
  assign nw04990 = ~(nw04989 | nw04982);
  assign nw04991 = nw04988 & ~(nw04990);
  assign nw05412[6] = nw04991 ^ nw04986;
  assign nw04992 = ~(\nr00016 [7] ^ \nr00017 [7]);
  assign nw05411[7] = ~nw04992;
  assign nw04993 = nw04991 | nw04986;
  assign nw04994 = nw04993 & ~(nw05413[6]);
  assign nw05412[7] = nw04994 ^ nw04992;
  assign nw04995 = ~(\nr00016 [8] ^ \nr00017 [8]);
  assign nw05411[8] = ~nw04995;
  assign nw04996 = nw05413[6] & ~(nw04992);
  assign nw04997 = nw04996 | nw05413[7];
  assign nw04998 = nw04992 | nw04986;
  assign nw04999 = ~(nw04998 | nw04988);
  assign nw05000 = nw04999 | nw04997;
  assign nw05001 = ~(nw04998 | nw04989);
  assign nw05002 = nw05001 & ~(nw04982);
  assign nw05003 = nw05002 | nw05000;
  assign nw05412[8] = nw05003 ^ nw05411[8];
  assign nw05004 = ~(\nr00016 [9] ^ \nr00017 [9]);
  assign nw05411[9] = ~nw05004;
  assign nw05005 = ~(nw05003 & nw05411[8]);
  assign nw05006 = nw05005 & ~(nw05413[8]);
  assign nw05412[9] = nw05006 ^ nw05004;
  assign nw05007 = ~(\nr00016 [10] ^ \nr00017 [10]);
  assign nw05411[10] = ~nw05007;
  assign nw05008 = nw05413[8] & ~(nw05004);
  assign nw05009 = ~(nw05008 | nw05413[9]);
  assign nw05010 = nw05004 | nw04995;
  assign nw05011 = nw05003 & ~(nw05010);
  assign nw05012 = nw05009 & ~(nw05011);
  assign nw05412[10] = nw05012 ^ nw05007;
  assign nw05013 = ~(\nr00016 [11] ^ \nr00017 [11]);
  assign nw05411[11] = ~nw05013;
  assign nw05014 = nw05012 | nw05007;
  assign nw05015 = nw05014 & ~(nw05413[10]);
  assign nw05412[11] = nw05015 ^ nw05013;
  assign nw05016 = ~(\nr00016 [12] ^ \nr00017 [12]);
  assign nw05411[12] = ~nw05016;
  assign nw05017 = nw05413[10] & ~(nw05013);
  assign nw05018 = nw05017 | nw05413[11];
  assign nw05019 = nw05013 | nw05007;
  assign nw05020 = ~(nw05019 | nw05009);
  assign nw05021 = nw05020 | nw05018;
  assign nw05022 = nw05019 | nw05010;
  assign nw05023 = nw05003 & ~(nw05022);
  assign nw05024 = ~(nw05023 | nw05021);
  assign nw05412[12] = nw05024 ^ nw05016;
  assign nw05025 = ~(\nr00016 [13] ^ \nr00017 [13]);
  assign nw05411[13] = ~nw05025;
  assign nw05026 = nw05411[12] & ~(nw05024);
  assign nw05027 = ~(nw05026 | nw05413[12]);
  assign nw05412[13] = nw05027 ^ nw05025;
  assign nw05028 = ~(\nr00016 [14] ^ \nr00017 [14]);
  assign nw05411[14] = ~nw05028;
  assign nw05029 = nw05413[12] & ~(nw05025);
  assign nw05030 = ~(nw05029 | nw05413[13]);
  assign nw05031 = nw05025 | nw05016;
  assign nw05032 = ~(nw05031 | nw05024);
  assign nw05033 = nw05030 & ~(nw05032);
  assign nw05412[14] = nw05033 ^ nw05028;
  assign nw05034 = ~(\nr00016 [15] ^ \nr00017 [15]);
  assign nw05411[15] = ~nw05034;
  assign nw05035 = nw05033 | nw05028;
  assign nw05036 = nw05035 & ~(nw05413[14]);
  assign nw05412[15] = nw05036 ^ nw05034;
  assign nw05037 = ~(\nr00016 [16] ^ \nr00017 [16]);
  assign nw05411[16] = ~nw05037;
  assign nw05038 = nw05413[14] & ~(nw05034);
  assign nw05039 = nw05038 | nw05413[15];
  assign nw05040 = nw05034 | nw05028;
  assign nw05041 = ~(nw05040 | nw05030);
  assign nw05042 = nw05041 | nw05039;
  assign nw05043 = nw05040 | nw05031;
  assign nw05044 = nw05021 & ~(nw05043);
  assign nw05045 = nw05044 | nw05042;
  assign nw05046 = nw05043 | nw05022;
  assign nw05047 = nw05003 & ~(nw05046);
  assign nw05048 = nw05047 | nw05045;
  assign nw05412[16] = nw05048 ^ nw05411[16];
  assign nw05049 = ~(\nr00016 [17] ^ \nr00017 [17]);
  assign nw05411[17] = ~nw05049;
  assign nw05050 = nw05048 & ~(nw05037);
  assign nw05051 = ~(nw05050 | nw05413[16]);
  assign nw05412[17] = nw05051 ^ nw05049;
  assign nw05052 = ~(\nr00016 [18] ^ \nr00017 [18]);
  assign nw05411[18] = ~nw05052;
  assign nw05053 = nw05413[16] & ~(nw05049);
  assign nw05054 = ~(nw05053 | nw05413[17]);
  assign nw05055 = nw05049 | nw05037;
  assign nw05056 = nw05048 & ~(nw05055);
  assign nw05057 = nw05054 & ~(nw05056);
  assign nw05412[18] = nw05057 ^ nw05052;
  assign nw05058 = ~(\nr00016 [19] ^ \nr00017 [19]);
  assign nw05411[19] = ~nw05058;
  assign nw05059 = nw05057 | nw05052;
  assign nw05060 = nw05059 & ~(nw05413[18]);
  assign nw05412[19] = nw05060 ^ nw05058;
  assign nw05061 = ~(\nr00016 [20] ^ \nr00017 [20]);
  assign nw05411[20] = ~nw05061;
  assign nw05062 = nw05413[18] & ~(nw05058);
  assign nw05063 = nw05062 | nw05413[19];
  assign nw05064 = nw05058 | nw05052;
  assign nw05065 = ~(nw05064 | nw05054);
  assign nw05066 = nw05065 | nw05063;
  assign nw05067 = nw05064 | nw05055;
  assign nw05068 = nw05048 & ~(nw05067);
  assign nw05069 = ~(nw05068 | nw05066);
  assign nw05412[20] = nw05069 ^ nw05061;
  assign nw05070 = ~(\nr00016 [21] ^ \nr00017 [21]);
  assign nw05411[21] = ~nw05070;
  assign nw05071 = nw05411[20] & ~(nw05069);
  assign nw05072 = ~(nw05071 | nw05413[20]);
  assign nw05412[21] = nw05072 ^ nw05070;
  assign nw05073 = ~(\nr00016 [22] ^ \nr00017 [22]);
  assign nw05411[22] = ~nw05073;
  assign nw05074 = nw05413[20] & ~(nw05070);
  assign nw05075 = ~(nw05074 | nw05413[21]);
  assign nw05076 = nw05070 | nw05061;
  assign nw05077 = ~(nw05076 | nw05069);
  assign nw05078 = nw05075 & ~(nw05077);
  assign nw05412[22] = nw05078 ^ nw05073;
  assign nw05079 = ~(\nr00016 [23] ^ \nr00017 [23]);
  assign nw05411[23] = ~nw05079;
  assign nw05080 = nw05078 | nw05073;
  assign nw05081 = nw05080 & ~(nw05413[22]);
  assign nw05412[23] = nw05081 ^ nw05079;
  assign nw05082 = ~(\nr00016 [24] ^ \nr00017 [24]);
  assign nw05411[24] = ~nw05082;
  assign nw05083 = nw05413[22] & ~(nw05079);
  assign nw05084 = ~(nw05083 | nw05413[23]);
  assign nw05085 = nw05079 | nw05073;
  assign nw05086 = ~(nw05085 | nw05075);
  assign nw05087 = nw05084 & ~(nw05086);
  assign nw05088 = nw05085 | nw05076;
  assign nw05089 = nw05066 & ~(nw05088);
  assign nw05090 = nw05087 & ~(nw05089);
  assign nw05091 = nw05088 | nw05067;
  assign nw05092 = nw05048 & ~(nw05091);
  assign nw05093 = nw05090 & ~(nw05092);
  assign nw05412[24] = nw05093 ^ nw05082;
  assign nw05094 = ~(\nr00016 [25] ^ \nr00017 [25]);
  assign nw05411[25] = ~nw05094;
  assign nw05095 = nw05411[24] & ~(nw05093);
  assign nw05096 = ~(nw05095 | nw05413[24]);
  assign nw05412[25] = nw05096 ^ nw05094;
  assign nw05097 = ~(\nr00016 [26] ^ \nr00017 [26]);
  assign nw05411[26] = ~nw05097;
  assign nw05098 = nw05413[24] & ~(nw05094);
  assign nw05099 = ~(nw05098 | nw05413[25]);
  assign nw05100 = nw05094 | nw05082;
  assign nw05101 = ~(nw05100 | nw05093);
  assign nw05102 = nw05099 & ~(nw05101);
  assign nw05412[26] = nw05102 ^ nw05097;
  assign nw05103 = ~(\nr00016 [27] ^ \nr00017 [27]);
  assign nw05411[27] = ~nw05103;
  assign nw05104 = nw05102 | nw05097;
  assign nw05105 = nw05104 & ~(nw05413[26]);
  assign nw05412[27] = nw05105 ^ nw05103;
  assign nw05106 = ~(\nr00016 [28] ^ \nr00017 [28]);
  assign nw05411[28] = ~nw05106;
  assign nw05107 = nw05413[26] & ~(nw05103);
  assign nw05108 = ~(nw05107 | nw05413[27]);
  assign nw05109 = nw05103 | nw05097;
  assign nw05110 = ~(nw05109 | nw05099);
  assign nw05111 = nw05108 & ~(nw05110);
  assign nw05112 = ~(nw05109 | nw05100);
  assign nw05113 = nw05112 & ~(nw05093);
  assign nw05114 = nw05111 & ~(nw05113);
  assign nw05412[28] = nw05114 ^ nw05106;
  assign nw05115 = ~(\nr00016 [29] ^ \nr00017 [29]);
  assign nw05411[29] = ~nw05115;
  assign nw05116 = nw05411[28] & ~(nw05114);
  assign nw05117 = ~(nw05116 | nw05413[28]);
  assign nw05412[29] = nw05117 ^ nw05115;
  assign nw05118 = ~(\nr00016 [30] ^ \nr00017 [30]);
  assign nw05411[30] = ~nw05118;
  assign nw05119 = nw05115 | ~(nw05413[28]);
  assign nw05120 = nw05119 & ~(nw05413[29]);
  assign nw05121 = nw05115 | nw05106;
  assign nw05122 = ~(nw05121 | nw05114);
  assign nw05123 = nw05120 & ~(nw05122);
  assign nw05412[30] = nw05123 ^ nw05118;
  assign nw05124 = ~(\nr00016 [31] ^ \nr00017 [31]);
  assign nw05411[31] = ~nw05124;
  assign nw05125 = nw05123 | nw05118;
  assign nw05126 = nw05125 & ~(nw05413[30]);
  assign nw05412[31] = nw05126 ^ nw05124;
  assign nw05411[0] = \nr00016 [0] ^ \nr00017 [0];
  assign nw05415[1] = \nw05427 [1] ^ \nw05427 [0];
  assign nw05127 = \nw05427 [1] & \nw05427 [0];
  assign nw05415[2] = nw05127 ^ \nw05427 [2];
  assign nw05128 = nw05127 & \nw05427 [2];
  assign nw05415[3] = nw05128 ^ \nw05427 [3];
  assign nw05129 = ~(\nw05427 [3] & \nw05427 [2]);
  assign nw05130 = nw05127 & ~(nw05129);
  assign nw05415[4] = nw05130 ^ \nw05427 [4];
  assign nw05131 = nw05130 & \nw05427 [4];
  assign nw05415[5] = nw05131 ^ \nw05427 [5];
  assign nw05132 = ~(\nw05427 [5] & \nw05427 [4]);
  assign nw05133 = nw05130 & ~(nw05132);
  assign nw05415[6] = nw05133 ^ \nw05427 [6];
  assign nw05134 = nw05133 & \nw05427 [6];
  assign nw05415[7] = nw05134 ^ \nw05427 [7];
  assign nw05135 = ~(\nw05427 [7] & \nw05427 [6]);
  assign nw05136 = nw05135 | nw05132;
  assign nw05137 = nw05130 & ~(nw05136);
  assign nw05415[8] = nw05137 ^ \nw05427 [8];
  assign nw05138 = nw05137 & \nw05427 [8];
  assign nw05415[9] = nw05138 ^ \nw05427 [9];
  assign nw05139 = ~(\nw05427 [9] & \nw05427 [8]);
  assign nw05140 = nw05137 & ~(nw05139);
  assign nw05415[10] = nw05140 ^ \nw05427 [10];
  assign nw05141 = nw05140 & \nw05427 [10];
  assign nw05415[11] = nw05141 ^ \nw05427 [11];
  assign nw05142 = ~(\nw05427 [11] & \nw05427 [10]);
  assign nw05143 = nw05142 | nw05139;
  assign nw05144 = nw05137 & ~(nw05143);
  assign nw05415[12] = nw05144 ^ \nw05427 [12];
  assign nw05145 = nw05144 & \nw05427 [12];
  assign nw05415[13] = nw05145 ^ \nw05427 [13];
  assign nw05146 = ~(\nw05427 [13] & \nw05427 [12]);
  assign nw05147 = nw05144 & ~(nw05146);
  assign nw05415[14] = nw05147 ^ \nw05427 [14];
  assign nw05148 = nw05147 & ~(nw04738);
  assign nw05415[15] = nw05148 ^ \nw05427 [15];
  assign nw05149 = nw05146 | nw04539;
  assign nw05150 = nw05149 | nw05143;
  assign nw05151 = nw05137 & ~(nw05150);
  assign nw05415[16] = nw05151 ^ \nw05427 [16];
  assign nw05152 = \nr00016 [0] & ~(\nr00017 [0]);
  assign nw05153 = nw05152 & ~(\nr00017 [1]);
  assign nw05154 = nw05153 & ~(\nr00017 [2]);
  assign nw05393 = nw05154 & ~(\nr00017 [3]);
  assign nw05155 = \nr00017 [0] ? \nr00016 [0] : \nr00016 [1];
  assign nw05156 = nw05155 & ~(\nr00017 [1]);
  assign nw05157 = nw05156 & ~(\nr00017 [2]);
  assign nw05394 = nw05157 & ~(\nr00017 [3]);
  assign nw05158 = \nr00017 [0] ? \nr00016 [1] : \nr00016 [2];
  assign nw05159 = \nr00017 [1] ? nw05152 : nw05158;
  assign nw05160 = nw05159 & ~(\nr00017 [2]);
  assign nw05395 = nw05160 & ~(\nr00017 [3]);
  assign nw05161 = \nr00017 [0] ? \nr00016 [2] : \nr00016 [3];
  assign nw05162 = \nr00017 [1] ? nw05155 : nw05161;
  assign nw05163 = nw05162 & ~(\nr00017 [2]);
  assign nw05396 = nw05163 & ~(\nr00017 [3]);
  assign nw05164 = \nr00017 [0] ? \nr00016 [3] : \nr00016 [4];
  assign nw05165 = \nr00017 [1] ? nw05158 : nw05164;
  assign nw05166 = \nr00017 [2] ? nw05153 : nw05165;
  assign nw05397 = nw05166 & ~(\nr00017 [3]);
  assign nw05167 = \nr00017 [0] ? \nr00016 [4] : \nr00016 [5];
  assign nw05168 = \nr00017 [1] ? nw05161 : nw05167;
  assign nw05169 = \nr00017 [2] ? nw05156 : nw05168;
  assign nw05398 = nw05169 & ~(\nr00017 [3]);
  assign nw05170 = \nr00017 [0] ? \nr00016 [5] : \nr00016 [6];
  assign nw05171 = \nr00017 [1] ? nw05164 : nw05170;
  assign nw05172 = \nr00017 [2] ? nw05159 : nw05171;
  assign nw05399 = nw05172 & ~(\nr00017 [3]);
  assign nw05173 = \nr00017 [0] ? \nr00016 [6] : \nr00016 [7];
  assign nw05174 = \nr00017 [1] ? nw05167 : nw05173;
  assign nw05175 = \nr00017 [2] ? nw05162 : nw05174;
  assign nw05400 = nw05175 & ~(\nr00017 [3]);
  assign nw05176 = \nr00017 [0] ? \nr00016 [7] : \nr00016 [8];
  assign nw05177 = \nr00017 [1] ? nw05170 : nw05176;
  assign nw05178 = \nr00017 [2] ? nw05165 : nw05177;
  assign nw05401 = \nr00017 [3] ? nw05154 : nw05178;
  assign nw05179 = \nr00017 [0] ? \nr00016 [8] : \nr00016 [9];
  assign nw05180 = \nr00017 [1] ? nw05173 : nw05179;
  assign nw05181 = \nr00017 [2] ? nw05168 : nw05180;
  assign nw05402 = \nr00017 [3] ? nw05157 : nw05181;
  assign nw05182 = \nr00017 [0] ? \nr00016 [9] : \nr00016 [10];
  assign nw05183 = \nr00017 [1] ? nw05176 : nw05182;
  assign nw05184 = \nr00017 [2] ? nw05171 : nw05183;
  assign nw05403 = \nr00017 [3] ? nw05160 : nw05184;
  assign nw05185 = \nr00017 [0] ? \nr00016 [10] : \nr00016 [11];
  assign nw05186 = \nr00017 [1] ? nw05179 : nw05185;
  assign nw05187 = \nr00017 [2] ? nw05174 : nw05186;
  assign nw05404 = \nr00017 [3] ? nw05163 : nw05187;
  assign nw05188 = \nr00017 [0] ? \nr00016 [11] : \nr00016 [12];
  assign nw05189 = \nr00017 [1] ? nw05182 : nw05188;
  assign nw05190 = \nr00017 [2] ? nw05177 : nw05189;
  assign nw05405 = \nr00017 [3] ? nw05166 : nw05190;
  assign nw05191 = \nr00017 [0] ? \nr00016 [12] : \nr00016 [13];
  assign nw05192 = \nr00017 [1] ? nw05185 : nw05191;
  assign nw05193 = \nr00017 [2] ? nw05180 : nw05192;
  assign nw05406 = \nr00017 [3] ? nw05169 : nw05193;
  assign nw05194 = \nr00017 [0] ? \nr00016 [13] : \nr00016 [14];
  assign nw05195 = \nr00017 [1] ? nw05188 : nw05194;
  assign nw05196 = \nr00017 [2] ? nw05183 : nw05195;
  assign nw05407 = \nr00017 [3] ? nw05172 : nw05196;
  assign nw05197 = \nr00017 [0] ? \nr00016 [14] : \nr00016 [15];
  assign nw05198 = \nr00017 [1] ? nw05191 : nw05197;
  assign nw05199 = \nr00017 [2] ? nw05186 : nw05198;
  assign nw05408 = \nr00017 [3] ? nw05175 : nw05199;
  assign nw05200 = \nr00017 [0] ? \nr00016 [15] : \nr00016 [16];
  assign nw05201 = \nr00017 [1] ? nw05194 : nw05200;
  assign nw05202 = \nr00017 [2] ? nw05189 : nw05201;
  assign nw05203 = \nr00017 [3] ? nw05178 : nw05202;
  assign nw05418[16] = \nr00017 [4] ? nw05393 : nw05203;
  assign nw05204 = \nr00017 [0] ? \nr00016 [16] : \nr00016 [17];
  assign nw05205 = \nr00017 [1] ? nw05197 : nw05204;
  assign nw05206 = \nr00017 [2] ? nw05192 : nw05205;
  assign nw05207 = \nr00017 [3] ? nw05181 : nw05206;
  assign nw05418[17] = \nr00017 [4] ? nw05394 : nw05207;
  assign nw05208 = \nr00017 [0] ? \nr00016 [17] : \nr00016 [18];
  assign nw05209 = \nr00017 [1] ? nw05200 : nw05208;
  assign nw05210 = \nr00017 [2] ? nw05195 : nw05209;
  assign nw05211 = \nr00017 [3] ? nw05184 : nw05210;
  assign nw05418[18] = \nr00017 [4] ? nw05395 : nw05211;
  assign nw05212 = \nr00017 [0] ? \nr00016 [18] : \nr00016 [19];
  assign nw05213 = \nr00017 [1] ? nw05204 : nw05212;
  assign nw05214 = \nr00017 [2] ? nw05198 : nw05213;
  assign nw05215 = \nr00017 [3] ? nw05187 : nw05214;
  assign nw05418[19] = \nr00017 [4] ? nw05396 : nw05215;
  assign nw05216 = \nr00017 [0] ? \nr00016 [19] : \nr00016 [20];
  assign nw05217 = \nr00017 [1] ? nw05208 : nw05216;
  assign nw05218 = \nr00017 [2] ? nw05201 : nw05217;
  assign nw05219 = \nr00017 [3] ? nw05190 : nw05218;
  assign nw05418[20] = \nr00017 [4] ? nw05397 : nw05219;
  assign nw05220 = \nr00017 [0] ? \nr00016 [20] : \nr00016 [21];
  assign nw05221 = \nr00017 [1] ? nw05212 : nw05220;
  assign nw05222 = \nr00017 [2] ? nw05205 : nw05221;
  assign nw05223 = \nr00017 [3] ? nw05193 : nw05222;
  assign nw05418[21] = \nr00017 [4] ? nw05398 : nw05223;
  assign nw05224 = \nr00017 [0] ? \nr00016 [21] : \nr00016 [22];
  assign nw05225 = \nr00017 [1] ? nw05216 : nw05224;
  assign nw05226 = \nr00017 [2] ? nw05209 : nw05225;
  assign nw05227 = \nr00017 [3] ? nw05196 : nw05226;
  assign nw05418[22] = \nr00017 [4] ? nw05399 : nw05227;
  assign nw05228 = \nr00017 [0] ? \nr00016 [22] : \nr00016 [23];
  assign nw05229 = \nr00017 [1] ? nw05220 : nw05228;
  assign nw05230 = \nr00017 [2] ? nw05213 : nw05229;
  assign nw05231 = \nr00017 [3] ? nw05199 : nw05230;
  assign nw05418[23] = \nr00017 [4] ? nw05400 : nw05231;
  assign nw05232 = \nr00017 [0] ? \nr00016 [23] : \nr00016 [24];
  assign nw05233 = \nr00017 [1] ? nw05224 : nw05232;
  assign nw05234 = \nr00017 [2] ? nw05217 : nw05233;
  assign nw05235 = \nr00017 [3] ? nw05202 : nw05234;
  assign nw05418[24] = \nr00017 [4] ? nw05401 : nw05235;
  assign nw05236 = \nr00017 [0] ? \nr00016 [24] : \nr00016 [25];
  assign nw05237 = \nr00017 [1] ? nw05228 : nw05236;
  assign nw05238 = \nr00017 [2] ? nw05221 : nw05237;
  assign nw05239 = \nr00017 [3] ? nw05206 : nw05238;
  assign nw05418[25] = \nr00017 [4] ? nw05402 : nw05239;
  assign nw05240 = \nr00017 [0] ? \nr00016 [25] : \nr00016 [26];
  assign nw05241 = \nr00017 [1] ? nw05232 : nw05240;
  assign nw05242 = \nr00017 [2] ? nw05225 : nw05241;
  assign nw05243 = \nr00017 [3] ? nw05210 : nw05242;
  assign nw05418[26] = \nr00017 [4] ? nw05403 : nw05243;
  assign nw05244 = \nr00017 [0] ? \nr00016 [26] : \nr00016 [27];
  assign nw05245 = \nr00017 [1] ? nw05236 : nw05244;
  assign nw05246 = \nr00017 [2] ? nw05229 : nw05245;
  assign nw05247 = \nr00017 [3] ? nw05214 : nw05246;
  assign nw05418[27] = \nr00017 [4] ? nw05404 : nw05247;
  assign nw05248 = \nr00017 [0] ? \nr00016 [27] : \nr00016 [28];
  assign nw05249 = \nr00017 [1] ? nw05240 : nw05248;
  assign nw05250 = \nr00017 [2] ? nw05233 : nw05249;
  assign nw05251 = \nr00017 [3] ? nw05218 : nw05250;
  assign nw05418[28] = \nr00017 [4] ? nw05405 : nw05251;
  assign nw05252 = \nr00017 [0] ? \nr00016 [28] : \nr00016 [29];
  assign nw05253 = \nr00017 [1] ? nw05244 : nw05252;
  assign nw05254 = \nr00017 [2] ? nw05237 : nw05253;
  assign nw05255 = \nr00017 [3] ? nw05222 : nw05254;
  assign nw05418[29] = \nr00017 [4] ? nw05406 : nw05255;
  assign nw05256 = \nr00017 [0] ? \nr00016 [29] : \nr00016 [30];
  assign nw05257 = \nr00017 [1] ? nw05248 : nw05256;
  assign nw05258 = \nr00017 [2] ? nw05241 : nw05257;
  assign nw05259 = \nr00017 [3] ? nw05226 : nw05258;
  assign nw05418[30] = \nr00017 [4] ? nw05407 : nw05259;
  assign nw05260 = \nr00017 [0] ? \nr00016 [30] : \nr00016 [31];
  assign nw05261 = \nr00017 [1] ? nw05252 : nw05260;
  assign nw05262 = \nr00017 [2] ? nw05245 : nw05261;
  assign nw05263 = \nr00017 [3] ? nw05230 : nw05262;
  assign nw05418[31] = \nr00017 [4] ? nw05408 : nw05263;
  assign nw05264 = \nr00017 [0] ? \nr00016 [1] : \nr00016 [0];
  assign nw05265 = \nr00017 [0] ? \nr00016 [3] : \nr00016 [2];
  assign nw05266 = \nr00017 [1] ? nw05265 : nw05264;
  assign nw05267 = \nr00017 [0] ? \nr00016 [5] : \nr00016 [4];
  assign nw05268 = \nr00017 [0] ? \nr00016 [7] : \nr00016 [6];
  assign nw05269 = \nr00017 [1] ? nw05268 : nw05267;
  assign nw05270 = \nr00017 [2] ? nw05269 : nw05266;
  assign nw05271 = \nr00017 [0] ? \nr00016 [9] : \nr00016 [8];
  assign nw05272 = \nr00017 [0] ? \nr00016 [11] : \nr00016 [10];
  assign nw05273 = \nr00017 [1] ? nw05272 : nw05271;
  assign nw05274 = \nr00017 [0] ? \nr00016 [13] : \nr00016 [12];
  assign nw05275 = \nr00017 [0] ? \nr00016 [15] : \nr00016 [14];
  assign nw05276 = \nr00017 [1] ? nw05275 : nw05274;
  assign nw05277 = \nr00017 [2] ? nw05276 : nw05273;
  assign nw05278 = \nr00017 [3] ? nw05277 : nw05270;
  assign nw05279 = \nr00017 [0] ? \nr00016 [17] : \nr00016 [16];
  assign nw05280 = \nr00017 [0] ? \nr00016 [19] : \nr00016 [18];
  assign nw05281 = \nr00017 [1] ? nw05280 : nw05279;
  assign nw05282 = \nr00017 [0] ? \nr00016 [21] : \nr00016 [20];
  assign nw05283 = \nr00017 [0] ? \nr00016 [23] : \nr00016 [22];
  assign nw05284 = \nr00017 [1] ? nw05283 : nw05282;
  assign nw05285 = \nr00017 [2] ? nw05284 : nw05281;
  assign nw05286 = \nr00017 [0] ? \nr00016 [25] : \nr00016 [24];
  assign nw05287 = \nr00017 [0] ? \nr00016 [27] : \nr00016 [26];
  assign nw05288 = \nr00017 [1] ? nw05287 : nw05286;
  assign nw05289 = \nr00017 [0] ? \nr00016 [29] : \nr00016 [28];
  assign nw05290 = \nr00017 [0] ? \nr00016 [31] : \nr00016 [30];
  assign nw05291 = \nr00017 [1] ? nw05290 : nw05289;
  assign nw05292 = \nr00017 [2] ? nw05291 : nw05288;
  assign nw05293 = \nr00017 [3] ? nw05292 : nw05285;
  assign nw05419[0] = \nr00017 [4] ? nw05293 : nw05278;
  assign nw05294 = \nr00017 [0] ? \nr00016 [2] : \nr00016 [1];
  assign nw05295 = \nr00017 [0] ? \nr00016 [4] : \nr00016 [3];
  assign nw05296 = \nr00017 [1] ? nw05295 : nw05294;
  assign nw05297 = \nr00017 [0] ? \nr00016 [6] : \nr00016 [5];
  assign nw05298 = \nr00017 [0] ? \nr00016 [8] : \nr00016 [7];
  assign nw05299 = \nr00017 [1] ? nw05298 : nw05297;
  assign nw05300 = \nr00017 [2] ? nw05299 : nw05296;
  assign nw05301 = \nr00017 [0] ? \nr00016 [10] : \nr00016 [9];
  assign nw05302 = \nr00017 [0] ? \nr00016 [12] : \nr00016 [11];
  assign nw05303 = \nr00017 [1] ? nw05302 : nw05301;
  assign nw05304 = \nr00017 [0] ? \nr00016 [14] : \nr00016 [13];
  assign nw05305 = \nr00017 [0] ? \nr00016 [16] : \nr00016 [15];
  assign nw05306 = \nr00017 [1] ? nw05305 : nw05304;
  assign nw05307 = \nr00017 [2] ? nw05306 : nw05303;
  assign nw05308 = \nr00017 [3] ? nw05307 : nw05300;
  assign nw05309 = \nr00017 [0] ? \nr00016 [18] : \nr00016 [17];
  assign nw05310 = \nr00017 [0] ? \nr00016 [20] : \nr00016 [19];
  assign nw05311 = \nr00017 [1] ? nw05310 : nw05309;
  assign nw05312 = \nr00017 [0] ? \nr00016 [22] : \nr00016 [21];
  assign nw05313 = \nr00017 [0] ? \nr00016 [24] : \nr00016 [23];
  assign nw05314 = \nr00017 [1] ? nw05313 : nw05312;
  assign nw05315 = \nr00017 [2] ? nw05314 : nw05311;
  assign nw05316 = \nr00017 [0] ? \nr00016 [26] : \nr00016 [25];
  assign nw05317 = \nr00017 [0] ? \nr00016 [28] : \nr00016 [27];
  assign nw05318 = \nr00017 [1] ? nw05317 : nw05316;
  assign nw05319 = \nr00017 [0] ? \nr00016 [30] : \nr00016 [29];
  assign nw05320 = \nr00016 [31] & ~(nw01373);
  assign nw05321 = \nr00017 [0] ? nw05320 : \nr00016 [31];
  assign nw05322 = \nr00017 [1] ? nw05321 : nw05319;
  assign nw05323 = \nr00017 [2] ? nw05322 : nw05318;
  assign nw05324 = \nr00017 [3] ? nw05323 : nw05315;
  assign nw05419[1] = \nr00017 [4] ? nw05324 : nw05308;
  assign nw05325 = \nr00017 [1] ? nw05267 : nw05265;
  assign nw05326 = \nr00017 [1] ? nw05271 : nw05268;
  assign nw05327 = \nr00017 [2] ? nw05326 : nw05325;
  assign nw05328 = \nr00017 [1] ? nw05274 : nw05272;
  assign nw05329 = \nr00017 [1] ? nw05279 : nw05275;
  assign nw05330 = \nr00017 [2] ? nw05329 : nw05328;
  assign nw05331 = \nr00017 [3] ? nw05330 : nw05327;
  assign nw05332 = \nr00017 [1] ? nw05282 : nw05280;
  assign nw05333 = \nr00017 [1] ? nw05286 : nw05283;
  assign nw05334 = \nr00017 [2] ? nw05333 : nw05332;
  assign nw05335 = \nr00017 [1] ? nw05289 : nw05287;
  assign nw05336 = \nr00017 [1] ? nw05320 : nw05290;
  assign nw05337 = \nr00017 [2] ? nw05336 : nw05335;
  assign nw05338 = \nr00017 [3] ? nw05337 : nw05334;
  assign nw05419[2] = \nr00017 [4] ? nw05338 : nw05331;
  assign nw05339 = \nr00017 [1] ? nw05297 : nw05295;
  assign nw05340 = \nr00017 [1] ? nw05301 : nw05298;
  assign nw05341 = \nr00017 [2] ? nw05340 : nw05339;
  assign nw05342 = \nr00017 [1] ? nw05304 : nw05302;
  assign nw05343 = \nr00017 [1] ? nw05309 : nw05305;
  assign nw05344 = \nr00017 [2] ? nw05343 : nw05342;
  assign nw05345 = \nr00017 [3] ? nw05344 : nw05341;
  assign nw05346 = \nr00017 [1] ? nw05312 : nw05310;
  assign nw05347 = \nr00017 [1] ? nw05316 : nw05313;
  assign nw05348 = \nr00017 [2] ? nw05347 : nw05346;
  assign nw05349 = \nr00017 [1] ? nw05319 : nw05317;
  assign nw05350 = \nr00017 [1] ? nw05320 : nw05321;
  assign nw05351 = \nr00017 [2] ? nw05350 : nw05349;
  assign nw05352 = \nr00017 [3] ? nw05351 : nw05348;
  assign nw05419[3] = \nr00017 [4] ? nw05352 : nw05345;
  assign nw05353 = \nr00017 [2] ? nw05273 : nw05269;
  assign nw05354 = \nr00017 [2] ? nw05281 : nw05276;
  assign nw05355 = \nr00017 [3] ? nw05354 : nw05353;
  assign nw05356 = \nr00017 [2] ? nw05288 : nw05284;
  assign nw05357 = \nr00017 [2] ? nw05320 : nw05291;
  assign nw05358 = \nr00017 [3] ? nw05357 : nw05356;
  assign nw05419[4] = \nr00017 [4] ? nw05358 : nw05355;
  assign nw05359 = \nr00017 [2] ? nw05303 : nw05299;
  assign nw05360 = \nr00017 [2] ? nw05311 : nw05306;
  assign nw05361 = \nr00017 [3] ? nw05360 : nw05359;
  assign nw05362 = \nr00017 [2] ? nw05318 : nw05314;
  assign nw05363 = \nr00017 [2] ? nw05320 : nw05322;
  assign nw05364 = \nr00017 [3] ? nw05363 : nw05362;
  assign nw05419[5] = \nr00017 [4] ? nw05364 : nw05361;
  assign nw05365 = \nr00017 [2] ? nw05328 : nw05326;
  assign nw05366 = \nr00017 [2] ? nw05332 : nw05329;
  assign nw05367 = \nr00017 [3] ? nw05366 : nw05365;
  assign nw05368 = \nr00017 [2] ? nw05335 : nw05333;
  assign nw05369 = \nr00017 [2] ? nw05320 : nw05336;
  assign nw05370 = \nr00017 [3] ? nw05369 : nw05368;
  assign nw05419[6] = \nr00017 [4] ? nw05370 : nw05367;
  assign nw05371 = \nr00017 [2] ? nw05342 : nw05340;
  assign nw05372 = \nr00017 [2] ? nw05346 : nw05343;
  assign nw05373 = \nr00017 [3] ? nw05372 : nw05371;
  assign nw05374 = \nr00017 [2] ? nw05349 : nw05347;
  assign nw05375 = \nr00017 [2] ? nw05320 : nw05350;
  assign nw05376 = \nr00017 [3] ? nw05375 : nw05374;
  assign nw05419[7] = \nr00017 [4] ? nw05376 : nw05373;
  assign nw05377 = \nr00017 [3] ? nw05285 : nw05277;
  assign nw05378 = \nr00017 [3] ? nw05320 : nw05292;
  assign nw05419[8] = \nr00017 [4] ? nw05378 : nw05377;
  assign nw05379 = \nr00017 [3] ? nw05315 : nw05307;
  assign nw05380 = \nr00017 [3] ? nw05320 : nw05323;
  assign nw05419[9] = \nr00017 [4] ? nw05380 : nw05379;
  assign nw05381 = \nr00017 [3] ? nw05334 : nw05330;
  assign nw05382 = \nr00017 [3] ? nw05320 : nw05337;
  assign nw05419[10] = \nr00017 [4] ? nw05382 : nw05381;
  assign nw05383 = \nr00017 [3] ? nw05348 : nw05344;
  assign nw05384 = \nr00017 [3] ? nw05320 : nw05351;
  assign nw05419[11] = \nr00017 [4] ? nw05384 : nw05383;
  assign nw05385 = \nr00017 [3] ? nw05356 : nw05354;
  assign nw05386 = \nr00017 [3] ? nw05320 : nw05357;
  assign nw05419[12] = \nr00017 [4] ? nw05386 : nw05385;
  assign nw05387 = \nr00017 [3] ? nw05362 : nw05360;
  assign nw05388 = \nr00017 [3] ? nw05320 : nw05363;
  assign nw05419[13] = \nr00017 [4] ? nw05388 : nw05387;
  assign nw05389 = \nr00017 [3] ? nw05368 : nw05366;
  assign nw05390 = \nr00017 [3] ? nw05320 : nw05369;
  assign nw05419[14] = \nr00017 [4] ? nw05390 : nw05389;
  assign nw05391 = \nr00017 [3] ? nw05374 : nw05372;
  assign nw05392 = \nr00017 [3] ? nw05320 : nw05375;
  assign nw05419[15] = \nr00017 [4] ? nw05392 : nw05391;
  assign nw05419[16] = \nr00017 [4] ? nw05320 : nw05293;
  assign nw05419[17] = \nr00017 [4] ? nw05320 : nw05324;
  assign nw05419[18] = \nr00017 [4] ? nw05320 : nw05338;
  assign nw05419[19] = \nr00017 [4] ? nw05320 : nw05352;
  assign nw05419[20] = \nr00017 [4] ? nw05320 : nw05358;
  assign nw05419[21] = \nr00017 [4] ? nw05320 : nw05364;
  assign nw05419[22] = \nr00017 [4] ? nw05320 : nw05370;
  assign nw05419[23] = \nr00017 [4] ? nw05320 : nw05376;
  assign nw05419[24] = \nr00017 [4] ? nw05320 : nw05378;
  assign nw05419[25] = \nr00017 [4] ? nw05320 : nw05380;
  assign nw05419[26] = \nr00017 [4] ? nw05320 : nw05382;
  assign nw05419[27] = \nr00017 [4] ? nw05320 : nw05384;
  assign nw05419[28] = \nr00017 [4] ? nw05320 : nw05386;
  assign nw05419[29] = \nr00017 [4] ? nw05320 : nw05388;
  assign nw05419[30] = \nr00017 [4] ? nw05320 : nw05390;
  assign nw05419[31] = \nr00017 [4] ? nw05320 : nw05392;
  always @(posedge clock_10_i)
    \nr00025 [0] <= nw00000;
  always @(posedge clock_10_i)
    \nr00025 [1] <= nw00001;
  always @(posedge clock_10_i)
    \nr00025 [2] <= nw00002;
  always @(posedge clock_10_i)
    \nr00025 [3] <= nw00003;
  always @(posedge clock_10_i)
    \nr00025 [4] <= nw00004;
  always @(posedge clock_10_i)
    \nr00025 [5] <= nw00005;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [0] <= 1'h0;
    else if (\nw05429 ) \nr00105 [0] <= ext_bus_data_o[0];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [1] <= 1'h0;
    else if (\nw05429 ) \nr00105 [1] <= ext_bus_data_o[1];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [2] <= 1'h0;
    else if (\nw05429 ) \nr00105 [2] <= ext_bus_data_o[2];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [3] <= 1'h0;
    else if (\nw05429 ) \nr00105 [3] <= ext_bus_data_o[3];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [4] <= 1'h0;
    else if (\nw05429 ) \nr00105 [4] <= ext_bus_data_o[4];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [5] <= 1'h0;
    else if (\nw05429 ) \nr00105 [5] <= ext_bus_data_o[5];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [6] <= 1'h0;
    else if (\nw05429 ) \nr00105 [6] <= ext_bus_data_o[6];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [7] <= 1'h0;
    else if (\nw05429 ) \nr00105 [7] <= ext_bus_data_o[7];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [8] <= 1'h0;
    else if (\nw05429 ) \nr00105 [8] <= ext_bus_data_o[8];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [9] <= 1'h0;
    else if (\nw05429 ) \nr00105 [9] <= ext_bus_data_o[9];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [10] <= 1'h0;
    else if (\nw05429 ) \nr00105 [10] <= ext_bus_data_o[10];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [11] <= 1'h0;
    else if (\nw05429 ) \nr00105 [11] <= ext_bus_data_o[11];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [12] <= 1'h0;
    else if (\nw05429 ) \nr00105 [12] <= ext_bus_data_o[12];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [13] <= 1'h0;
    else if (\nw05429 ) \nr00105 [13] <= ext_bus_data_o[13];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [14] <= 1'h0;
    else if (\nw05429 ) \nr00105 [14] <= ext_bus_data_o[14];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [15] <= 1'h0;
    else if (\nw05429 ) \nr00105 [15] <= ext_bus_data_o[15];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [16] <= 1'h0;
    else if (\nw05429 ) \nr00105 [16] <= ext_bus_data_o[16];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [17] <= 1'h0;
    else if (\nw05429 ) \nr00105 [17] <= ext_bus_data_o[17];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [18] <= 1'h0;
    else if (\nw05429 ) \nr00105 [18] <= ext_bus_data_o[18];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [19] <= 1'h0;
    else if (\nw05429 ) \nr00105 [19] <= ext_bus_data_o[19];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [20] <= 1'h0;
    else if (\nw05429 ) \nr00105 [20] <= ext_bus_data_o[20];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [21] <= 1'h0;
    else if (\nw05429 ) \nr00105 [21] <= ext_bus_data_o[21];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [22] <= 1'h0;
    else if (\nw05429 ) \nr00105 [22] <= ext_bus_data_o[22];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [23] <= 1'h0;
    else if (\nw05429 ) \nr00105 [23] <= ext_bus_data_o[23];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [24] <= 1'h0;
    else if (\nw05429 ) \nr00105 [24] <= ext_bus_data_o[24];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [25] <= 1'h0;
    else if (\nw05429 ) \nr00105 [25] <= ext_bus_data_o[25];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [26] <= 1'h0;
    else if (\nw05429 ) \nr00105 [26] <= ext_bus_data_o[26];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [27] <= 1'h0;
    else if (\nw05429 ) \nr00105 [27] <= ext_bus_data_o[27];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [28] <= 1'h0;
    else if (\nw05429 ) \nr00105 [28] <= ext_bus_data_o[28];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [29] <= 1'h0;
    else if (\nw05429 ) \nr00105 [29] <= ext_bus_data_o[29];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [30] <= 1'h0;
    else if (\nw05429 ) \nr00105 [30] <= ext_bus_data_o[30];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00105 [31] <= 1'h0;
    else if (\nw05429 ) \nr00105 [31] <= ext_bus_data_o[31];
  reg \nr00106[0]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[0]  <= 1'h0;
    else \nr00106[0]  <= nw05414[0];
  assign \nw05427 [0] = \nr00106[0] ;
  reg \nr00106[1]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[1]  <= 1'h0;
    else \nr00106[1]  <= nw05415[1];
  assign \nw05427 [1] = \nr00106[1] ;
  reg \nr00106[2]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[2]  <= 1'h0;
    else \nr00106[2]  <= nw05415[2];
  assign \nw05427 [2] = \nr00106[2] ;
  reg \nr00106[3]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[3]  <= 1'h0;
    else \nr00106[3]  <= nw05415[3];
  assign \nw05427 [3] = \nr00106[3] ;
  reg \nr00106[4]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[4]  <= 1'h0;
    else \nr00106[4]  <= nw05415[4];
  assign \nw05427 [4] = \nr00106[4] ;
  reg \nr00106[5]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[5]  <= 1'h0;
    else \nr00106[5]  <= nw05415[5];
  assign \nw05427 [5] = \nr00106[5] ;
  reg \nr00106[6]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[6]  <= 1'h0;
    else \nr00106[6]  <= nw05415[6];
  assign \nw05427 [6] = \nr00106[6] ;
  reg \nr00106[7]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[7]  <= 1'h0;
    else \nr00106[7]  <= nw05415[7];
  assign \nw05427 [7] = \nr00106[7] ;
  reg \nr00106[8]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[8]  <= 1'h0;
    else \nr00106[8]  <= nw05415[8];
  assign \nw05427 [8] = \nr00106[8] ;
  reg \nr00106[9]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[9]  <= 1'h0;
    else \nr00106[9]  <= nw05415[9];
  assign \nw05427 [9] = \nr00106[9] ;
  reg \nr00106[10]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[10]  <= 1'h0;
    else \nr00106[10]  <= nw05415[10];
  assign \nw05427 [10] = \nr00106[10] ;
  reg \nr00106[11]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[11]  <= 1'h0;
    else \nr00106[11]  <= nw05415[11];
  assign \nw05427 [11] = \nr00106[11] ;
  reg \nr00106[12]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[12]  <= 1'h0;
    else \nr00106[12]  <= nw05415[12];
  assign \nw05427 [12] = \nr00106[12] ;
  reg \nr00106[13]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[13]  <= 1'h0;
    else \nr00106[13]  <= nw05415[13];
  assign \nw05427 [13] = \nr00106[13] ;
  reg \nr00106[14]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[14]  <= 1'h0;
    else \nr00106[14]  <= nw05415[14];
  assign \nw05427 [14] = \nr00106[14] ;
  reg \nr00106[15]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[15]  <= 1'h0;
    else \nr00106[15]  <= nw05415[15];
  assign \nw05427 [15] = \nr00106[15] ;
  reg \nr00106[16]  = 1'h0;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00106[16]  <= 1'h0;
    else \nr00106[16]  <= nw05415[16];
  assign \nw05427 [16] = \nr00106[16] ;
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[0] <= 1'h0;
    else if (nw00040) nr00009[0] <= nw05421[0];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[1] <= 1'h0;
    else if (nw00040) nr00009[1] <= nw05421[1];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[2] <= 1'h0;
    else if (nw00040) nr00009[2] <= nw05421[2];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[3] <= 1'h0;
    else if (nw00040) nr00009[3] <= nw05421[3];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[4] <= 1'h0;
    else if (nw00040) nr00009[4] <= nw05421[4];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[5] <= 1'h0;
    else if (nw00040) nr00009[5] <= nw05421[5];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[6] <= 1'h0;
    else if (nw00040) nr00009[6] <= nw05421[6];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[7] <= 1'h0;
    else if (nw00040) nr00009[7] <= nw05421[7];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[8] <= 1'h0;
    else if (nw00040) nr00009[8] <= nw05421[8];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[9] <= 1'h0;
    else if (nw00040) nr00009[9] <= nw05421[9];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[10] <= 1'h0;
    else if (nw00040) nr00009[10] <= nw05421[10];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[11] <= 1'h0;
    else if (nw00040) nr00009[11] <= nw05421[11];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[12] <= 1'h0;
    else if (nw00040) nr00009[12] <= nw05421[12];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[13] <= 1'h0;
    else if (nw00040) nr00009[13] <= nw05421[13];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[14] <= 1'h0;
    else if (nw00040) nr00009[14] <= nw05421[14];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[15] <= 1'h0;
    else if (nw00040) nr00009[15] <= nw05421[15];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[16] <= 1'h0;
    else if (nw00040) nr00009[16] <= nw05421[16];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[17] <= 1'h0;
    else if (nw00040) nr00009[17] <= nw05421[17];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[18] <= 1'h0;
    else if (nw00040) nr00009[18] <= nw05421[18];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[19] <= 1'h0;
    else if (nw00040) nr00009[19] <= nw05421[19];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[20] <= 1'h0;
    else if (nw00040) nr00009[20] <= nw05421[20];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[21] <= 1'h0;
    else if (nw00040) nr00009[21] <= nw05421[21];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[22] <= 1'h0;
    else if (nw00040) nr00009[22] <= nw05421[22];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[23] <= 1'h0;
    else if (nw00040) nr00009[23] <= nw05421[23];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[24] <= 1'h0;
    else if (nw00040) nr00009[24] <= nw05421[24];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[25] <= 1'h0;
    else if (nw00040) nr00009[25] <= nw05421[25];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[26] <= 1'h0;
    else if (nw00040) nr00009[26] <= nw05421[26];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[27] <= 1'h0;
    else if (nw00040) nr00009[27] <= nw05421[27];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[28] <= 1'h0;
    else if (nw00040) nr00009[28] <= nw05421[28];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[29] <= 1'h0;
    else if (nw00040) nr00009[29] <= nw05421[29];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[30] <= 1'h0;
    else if (nw00040) nr00009[30] <= nw05421[30];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) nr00009[31] <= 1'h0;
    else if (nw00040) nr00009[31] <= nw05421[31];
  always @(posedge clock_10_i)
    \nr00103 [0] <= nw05420[0];
  always @(posedge clock_10_i)
    \nr00103 [1] <= nw05420[1];
  always @(posedge clock_10_i)
    \nr00103 [2] <= nw05420[2];
  always @(posedge clock_10_i)
    \nr00103 [3] <= nw05420[3];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [0] <= 1'h0;
    else if (\nw05428 ) \nr00104 [0] <= ext_bus_data_o[0];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [1] <= 1'h0;
    else if (\nw05428 ) \nr00104 [1] <= ext_bus_data_o[1];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [2] <= 1'h0;
    else if (\nw05428 ) \nr00104 [2] <= ext_bus_data_o[2];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [3] <= 1'h0;
    else if (\nw05428 ) \nr00104 [3] <= ext_bus_data_o[3];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [4] <= 1'h0;
    else if (\nw05428 ) \nr00104 [4] <= ext_bus_data_o[4];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [5] <= 1'h0;
    else if (\nw05428 ) \nr00104 [5] <= ext_bus_data_o[5];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [6] <= 1'h0;
    else if (\nw05428 ) \nr00104 [6] <= ext_bus_data_o[6];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [7] <= 1'h0;
    else if (\nw05428 ) \nr00104 [7] <= ext_bus_data_o[7];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [8] <= 1'h0;
    else if (\nw05428 ) \nr00104 [8] <= ext_bus_data_o[8];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [9] <= 1'h0;
    else if (\nw05428 ) \nr00104 [9] <= ext_bus_data_o[9];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [10] <= 1'h0;
    else if (\nw05428 ) \nr00104 [10] <= ext_bus_data_o[10];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [11] <= 1'h0;
    else if (\nw05428 ) \nr00104 [11] <= ext_bus_data_o[11];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [12] <= 1'h0;
    else if (\nw05428 ) \nr00104 [12] <= ext_bus_data_o[12];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [13] <= 1'h0;
    else if (\nw05428 ) \nr00104 [13] <= ext_bus_data_o[13];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [14] <= 1'h0;
    else if (\nw05428 ) \nr00104 [14] <= ext_bus_data_o[14];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [15] <= 1'h0;
    else if (\nw05428 ) \nr00104 [15] <= ext_bus_data_o[15];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [16] <= 1'h0;
    else if (\nw05428 ) \nr00104 [16] <= ext_bus_data_o[16];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [17] <= 1'h0;
    else if (\nw05428 ) \nr00104 [17] <= ext_bus_data_o[17];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [18] <= 1'h0;
    else if (\nw05428 ) \nr00104 [18] <= ext_bus_data_o[18];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [19] <= 1'h0;
    else if (\nw05428 ) \nr00104 [19] <= ext_bus_data_o[19];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [20] <= 1'h0;
    else if (\nw05428 ) \nr00104 [20] <= ext_bus_data_o[20];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [21] <= 1'h0;
    else if (\nw05428 ) \nr00104 [21] <= ext_bus_data_o[21];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [22] <= 1'h0;
    else if (\nw05428 ) \nr00104 [22] <= ext_bus_data_o[22];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [23] <= 1'h0;
    else if (\nw05428 ) \nr00104 [23] <= ext_bus_data_o[23];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [24] <= 1'h0;
    else if (\nw05428 ) \nr00104 [24] <= ext_bus_data_o[24];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [25] <= 1'h0;
    else if (\nw05428 ) \nr00104 [25] <= ext_bus_data_o[25];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [26] <= 1'h0;
    else if (\nw05428 ) \nr00104 [26] <= ext_bus_data_o[26];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [27] <= 1'h0;
    else if (\nw05428 ) \nr00104 [27] <= ext_bus_data_o[27];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [28] <= 1'h0;
    else if (\nw05428 ) \nr00104 [28] <= ext_bus_data_o[28];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [29] <= 1'h0;
    else if (\nw05428 ) \nr00104 [29] <= ext_bus_data_o[29];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [30] <= 1'h0;
    else if (\nw05428 ) \nr00104 [30] <= ext_bus_data_o[30];
  always @(posedge clock_10_i)
    if (reset_effectivo_o) \nr00104 [31] <= 1'h0;
    else if (\nw05428 ) \nr00104 [31] <= ext_bus_data_o[31];
  always @(posedge clock_10_i)
    \nr00007 [0] <= \nr00006 [0];
  always @(posedge clock_10_i)
    \nr00007 [1] <= \nr00006 [1];
  always @(posedge clock_10_i)
    \nr00007 [2] <= \nr00006 [2];
  always @(posedge clock_10_i)
    \nr00007 [3] <= \nr00006 [3];
  always @(posedge clock_10_i)
    \nr00007 [4] <= \nr00006 [4];
  always @(posedge clock_10_i)
    \nr00007 [5] <= \nr00006 [5];
  always @(posedge clock_10_i)
    \nr00007 [6] <= \nr00006 [6];
  always @(posedge clock_10_i)
    \nr00007 [7] <= \nr00006 [7];
  always @(posedge clock_10_i)
    \nr00007 [8] <= \nr00006 [8];
  always @(posedge clock_10_i)
    \nr00007 [9] <= \nr00006 [9];
  always @(posedge clock_10_i)
    \nr00007 [10] <= \nr00006 [10];
  always @(posedge clock_10_i)
    \nr00007 [11] <= \nr00006 [11];
  always @(posedge clock_10_i)
    \nr00007 [12] <= \nr00006 [12];
  always @(posedge clock_10_i)
    \nr00007 [13] <= \nr00006 [13];
  always @(posedge clock_10_i)
    \nr00007 [14] <= \nr00006 [14];
  always @(posedge clock_10_i)
    \nr00007 [15] <= \nr00006 [15];
  always @(posedge clock_10_i)
    \nr00006 [0] <= \nr00005 [0];
  always @(posedge clock_10_i)
    \nr00006 [1] <= \nr00005 [1];
  always @(posedge clock_10_i)
    \nr00006 [2] <= \nr00005 [2];
  always @(posedge clock_10_i)
    \nr00006 [3] <= \nr00005 [3];
  always @(posedge clock_10_i)
    \nr00006 [4] <= \nr00005 [4];
  always @(posedge clock_10_i)
    \nr00006 [5] <= \nr00005 [5];
  always @(posedge clock_10_i)
    \nr00006 [6] <= \nr00005 [6];
  always @(posedge clock_10_i)
    \nr00006 [7] <= \nr00005 [7];
  always @(posedge clock_10_i)
    \nr00006 [8] <= \nr00005 [8];
  always @(posedge clock_10_i)
    \nr00006 [9] <= \nr00005 [9];
  always @(posedge clock_10_i)
    \nr00006 [10] <= \nr00005 [10];
  always @(posedge clock_10_i)
    \nr00006 [11] <= \nr00005 [11];
  always @(posedge clock_10_i)
    \nr00006 [12] <= \nr00005 [12];
  always @(posedge clock_10_i)
    \nr00006 [13] <= \nr00005 [13];
  always @(posedge clock_10_i)
    \nr00006 [14] <= \nr00005 [14];
  always @(posedge clock_10_i)
    \nr00006 [15] <= \nr00005 [15];
  always @(posedge clock_10_i)
    \nr00005 [0] <= sw_i[0];
  always @(posedge clock_10_i)
    \nr00005 [1] <= sw_i[1];
  always @(posedge clock_10_i)
    \nr00005 [2] <= sw_i[2];
  always @(posedge clock_10_i)
    \nr00005 [3] <= sw_i[3];
  always @(posedge clock_10_i)
    \nr00005 [4] <= sw_i[4];
  always @(posedge clock_10_i)
    \nr00005 [5] <= sw_i[5];
  always @(posedge clock_10_i)
    \nr00005 [6] <= sw_i[6];
  always @(posedge clock_10_i)
    \nr00005 [7] <= sw_i[7];
  always @(posedge clock_10_i)
    \nr00005 [8] <= sw_i[8];
  always @(posedge clock_10_i)
    \nr00005 [9] <= sw_i[9];
  always @(posedge clock_10_i)
    \nr00005 [10] <= sw_i[10];
  always @(posedge clock_10_i)
    \nr00005 [11] <= sw_i[11];
  always @(posedge clock_10_i)
    \nr00005 [12] <= sw_i[12];
  always @(posedge clock_10_i)
    \nr00005 [13] <= sw_i[13];
  always @(posedge clock_10_i)
    \nr00005 [14] <= sw_i[14];
  always @(posedge clock_10_i)
    \nr00005 [15] <= sw_i[15];
  always @(posedge clock_10_i)
    \nr00004 [0] <= \nr00003 [0];
  always @(posedge clock_10_i)
    \nr00004 [1] <= \nr00003 [1];
  always @(posedge clock_10_i)
    \nr00004 [2] <= \nr00003 [2];
  always @(posedge clock_10_i)
    \nr00004 [3] <= \nr00003 [3];
  always @(posedge clock_10_i)
    \nr00003 [0] <= \nr00002 [0];
  always @(posedge clock_10_i)
    \nr00003 [1] <= \nr00002 [1];
  always @(posedge clock_10_i)
    \nr00003 [2] <= \nr00002 [2];
  always @(posedge clock_10_i)
    \nr00003 [3] <= \nr00002 [3];
  always @(posedge clock_10_i)
    \nr00002 [0] <= btn_i[0];
  always @(posedge clock_10_i)
    \nr00002 [1] <= btn_i[1];
  always @(posedge clock_10_i)
    \nr00002 [2] <= btn_i[2];
  always @(posedge clock_10_i)
    \nr00002 [3] <= btn_i[3];
  always @(posedge clock_10_i)
    if (nw00042) \nr00017 [0] <= nw00097;
  always @(posedge clock_10_i)
    if (nw00042) \nr00017 [1] <= nw00098;
  always @(posedge clock_10_i)
    if (nw00042) \nr00017 [2] <= nw00099;
  always @(posedge clock_10_i)
    if (nw00042) \nr00017 [3] <= nw00100;
  always @(posedge clock_10_i)
    if (nw00042) \nr00017 [4] <= nw00101;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [0] <= 1'h0;
      else \nr00071[30] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [1] <= 1'h0;
      else \nr00071[30] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [2] <= 1'h0;
      else \nr00071[30] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [3] <= 1'h0;
      else \nr00071[30] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [4] <= 1'h0;
      else \nr00071[30] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [5] <= 1'h0;
      else \nr00071[30] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [6] <= 1'h0;
      else \nr00071[30] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [7] <= 1'h0;
      else \nr00071[30] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [8] <= 1'h0;
      else \nr00071[30] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [9] <= 1'h0;
      else \nr00071[30] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [10] <= 1'h0;
      else \nr00071[30] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [11] <= 1'h0;
      else \nr00071[30] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [12] <= 1'h0;
      else \nr00071[30] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [13] <= 1'h0;
      else \nr00071[30] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [14] <= 1'h0;
      else \nr00071[30] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [15] <= 1'h0;
      else \nr00071[30] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [16] <= 1'h0;
      else \nr00071[30] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [17] <= 1'h0;
      else \nr00071[30] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [18] <= 1'h0;
      else \nr00071[30] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [19] <= 1'h0;
      else \nr00071[30] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [20] <= 1'h0;
      else \nr00071[30] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [21] <= 1'h0;
      else \nr00071[30] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [22] <= 1'h0;
      else \nr00071[30] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [23] <= 1'h0;
      else \nr00071[30] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [24] <= 1'h0;
      else \nr00071[30] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [25] <= 1'h0;
      else \nr00071[30] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [26] <= 1'h0;
      else \nr00071[30] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [27] <= 1'h0;
      else \nr00071[30] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [28] <= 1'h0;
      else \nr00071[30] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [29] <= 1'h0;
      else \nr00071[30] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [30] <= 1'h0;
      else \nr00071[30] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00017)
      if (!nw00407) \nr00071[30] [31] <= 1'h0;
      else \nr00071[30] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [0] <= 1'h0;
      else \nr00071[29] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [1] <= 1'h0;
      else \nr00071[29] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [2] <= 1'h0;
      else \nr00071[29] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [3] <= 1'h0;
      else \nr00071[29] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [4] <= 1'h0;
      else \nr00071[29] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [5] <= 1'h0;
      else \nr00071[29] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [6] <= 1'h0;
      else \nr00071[29] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [7] <= 1'h0;
      else \nr00071[29] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [8] <= 1'h0;
      else \nr00071[29] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [9] <= 1'h0;
      else \nr00071[29] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [10] <= 1'h0;
      else \nr00071[29] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [11] <= 1'h0;
      else \nr00071[29] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [12] <= 1'h0;
      else \nr00071[29] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [13] <= 1'h0;
      else \nr00071[29] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [14] <= 1'h0;
      else \nr00071[29] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [15] <= 1'h0;
      else \nr00071[29] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [16] <= 1'h0;
      else \nr00071[29] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [17] <= 1'h0;
      else \nr00071[29] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [18] <= 1'h0;
      else \nr00071[29] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [19] <= 1'h0;
      else \nr00071[29] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [20] <= 1'h0;
      else \nr00071[29] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [21] <= 1'h0;
      else \nr00071[29] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [22] <= 1'h0;
      else \nr00071[29] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [23] <= 1'h0;
      else \nr00071[29] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [24] <= 1'h0;
      else \nr00071[29] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [25] <= 1'h0;
      else \nr00071[29] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [26] <= 1'h0;
      else \nr00071[29] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [27] <= 1'h0;
      else \nr00071[29] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [28] <= 1'h0;
      else \nr00071[29] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [29] <= 1'h0;
      else \nr00071[29] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [30] <= 1'h0;
      else \nr00071[29] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00019)
      if (!nw00405) \nr00071[29] [31] <= 1'h0;
      else \nr00071[29] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [0] <= 1'h0;
      else \nr00071[28] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [1] <= 1'h0;
      else \nr00071[28] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [2] <= 1'h0;
      else \nr00071[28] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [3] <= 1'h0;
      else \nr00071[28] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [4] <= 1'h0;
      else \nr00071[28] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [5] <= 1'h0;
      else \nr00071[28] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [6] <= 1'h0;
      else \nr00071[28] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [7] <= 1'h0;
      else \nr00071[28] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [8] <= 1'h0;
      else \nr00071[28] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [9] <= 1'h0;
      else \nr00071[28] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [10] <= 1'h0;
      else \nr00071[28] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [11] <= 1'h0;
      else \nr00071[28] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [12] <= 1'h0;
      else \nr00071[28] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [13] <= 1'h0;
      else \nr00071[28] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [14] <= 1'h0;
      else \nr00071[28] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [15] <= 1'h0;
      else \nr00071[28] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [16] <= 1'h0;
      else \nr00071[28] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [17] <= 1'h0;
      else \nr00071[28] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [18] <= 1'h0;
      else \nr00071[28] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [19] <= 1'h0;
      else \nr00071[28] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [20] <= 1'h0;
      else \nr00071[28] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [21] <= 1'h0;
      else \nr00071[28] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [22] <= 1'h0;
      else \nr00071[28] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [23] <= 1'h0;
      else \nr00071[28] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [24] <= 1'h0;
      else \nr00071[28] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [25] <= 1'h0;
      else \nr00071[28] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [26] <= 1'h0;
      else \nr00071[28] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [27] <= 1'h0;
      else \nr00071[28] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [28] <= 1'h0;
      else \nr00071[28] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [29] <= 1'h0;
      else \nr00071[28] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [30] <= 1'h0;
      else \nr00071[28] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00020)
      if (!nw00404) \nr00071[28] [31] <= 1'h0;
      else \nr00071[28] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [0] <= 1'h0;
      else \nr00071[27] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [1] <= 1'h0;
      else \nr00071[27] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [2] <= 1'h0;
      else \nr00071[27] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [3] <= 1'h0;
      else \nr00071[27] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [4] <= 1'h0;
      else \nr00071[27] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [5] <= 1'h0;
      else \nr00071[27] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [6] <= 1'h0;
      else \nr00071[27] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [7] <= 1'h0;
      else \nr00071[27] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [8] <= 1'h0;
      else \nr00071[27] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [9] <= 1'h0;
      else \nr00071[27] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [10] <= 1'h0;
      else \nr00071[27] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [11] <= 1'h0;
      else \nr00071[27] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [12] <= 1'h0;
      else \nr00071[27] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [13] <= 1'h0;
      else \nr00071[27] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [14] <= 1'h0;
      else \nr00071[27] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [15] <= 1'h0;
      else \nr00071[27] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [16] <= 1'h0;
      else \nr00071[27] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [17] <= 1'h0;
      else \nr00071[27] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [18] <= 1'h0;
      else \nr00071[27] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [19] <= 1'h0;
      else \nr00071[27] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [20] <= 1'h0;
      else \nr00071[27] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [21] <= 1'h0;
      else \nr00071[27] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [22] <= 1'h0;
      else \nr00071[27] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [23] <= 1'h0;
      else \nr00071[27] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [24] <= 1'h0;
      else \nr00071[27] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [25] <= 1'h0;
      else \nr00071[27] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [26] <= 1'h0;
      else \nr00071[27] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [27] <= 1'h0;
      else \nr00071[27] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [28] <= 1'h0;
      else \nr00071[27] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [29] <= 1'h0;
      else \nr00071[27] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [30] <= 1'h0;
      else \nr00071[27] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00021)
      if (!nw00403) \nr00071[27] [31] <= 1'h0;
      else \nr00071[27] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [0] <= 1'h0;
      else \nr00071[26] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [1] <= 1'h0;
      else \nr00071[26] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [2] <= 1'h0;
      else \nr00071[26] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [3] <= 1'h0;
      else \nr00071[26] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [4] <= 1'h0;
      else \nr00071[26] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [5] <= 1'h0;
      else \nr00071[26] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [6] <= 1'h0;
      else \nr00071[26] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [7] <= 1'h0;
      else \nr00071[26] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [8] <= 1'h0;
      else \nr00071[26] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [9] <= 1'h0;
      else \nr00071[26] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [10] <= 1'h0;
      else \nr00071[26] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [11] <= 1'h0;
      else \nr00071[26] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [12] <= 1'h0;
      else \nr00071[26] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [13] <= 1'h0;
      else \nr00071[26] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [14] <= 1'h0;
      else \nr00071[26] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [15] <= 1'h0;
      else \nr00071[26] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [16] <= 1'h0;
      else \nr00071[26] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [17] <= 1'h0;
      else \nr00071[26] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [18] <= 1'h0;
      else \nr00071[26] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [19] <= 1'h0;
      else \nr00071[26] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [20] <= 1'h0;
      else \nr00071[26] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [21] <= 1'h0;
      else \nr00071[26] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [22] <= 1'h0;
      else \nr00071[26] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [23] <= 1'h0;
      else \nr00071[26] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [24] <= 1'h0;
      else \nr00071[26] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [25] <= 1'h0;
      else \nr00071[26] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [26] <= 1'h0;
      else \nr00071[26] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [27] <= 1'h0;
      else \nr00071[26] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [28] <= 1'h0;
      else \nr00071[26] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [29] <= 1'h0;
      else \nr00071[26] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [30] <= 1'h0;
      else \nr00071[26] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00022)
      if (!nw00402) \nr00071[26] [31] <= 1'h0;
      else \nr00071[26] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [0] <= 1'h0;
      else \nr00071[25] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [1] <= 1'h0;
      else \nr00071[25] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [2] <= 1'h0;
      else \nr00071[25] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [3] <= 1'h0;
      else \nr00071[25] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [4] <= 1'h0;
      else \nr00071[25] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [5] <= 1'h0;
      else \nr00071[25] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [6] <= 1'h0;
      else \nr00071[25] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [7] <= 1'h0;
      else \nr00071[25] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [8] <= 1'h0;
      else \nr00071[25] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [9] <= 1'h0;
      else \nr00071[25] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [10] <= 1'h0;
      else \nr00071[25] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [11] <= 1'h0;
      else \nr00071[25] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [12] <= 1'h0;
      else \nr00071[25] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [13] <= 1'h0;
      else \nr00071[25] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [14] <= 1'h0;
      else \nr00071[25] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [15] <= 1'h0;
      else \nr00071[25] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [16] <= 1'h0;
      else \nr00071[25] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [17] <= 1'h0;
      else \nr00071[25] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [18] <= 1'h0;
      else \nr00071[25] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [19] <= 1'h0;
      else \nr00071[25] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [20] <= 1'h0;
      else \nr00071[25] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [21] <= 1'h0;
      else \nr00071[25] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [22] <= 1'h0;
      else \nr00071[25] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [23] <= 1'h0;
      else \nr00071[25] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [24] <= 1'h0;
      else \nr00071[25] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [25] <= 1'h0;
      else \nr00071[25] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [26] <= 1'h0;
      else \nr00071[25] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [27] <= 1'h0;
      else \nr00071[25] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [28] <= 1'h0;
      else \nr00071[25] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [29] <= 1'h0;
      else \nr00071[25] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [30] <= 1'h0;
      else \nr00071[25] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00023)
      if (!nw00401) \nr00071[25] [31] <= 1'h0;
      else \nr00071[25] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [0] <= 1'h0;
      else \nr00071[24] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [1] <= 1'h0;
      else \nr00071[24] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [2] <= 1'h0;
      else \nr00071[24] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [3] <= 1'h0;
      else \nr00071[24] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [4] <= 1'h0;
      else \nr00071[24] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [5] <= 1'h0;
      else \nr00071[24] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [6] <= 1'h0;
      else \nr00071[24] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [7] <= 1'h0;
      else \nr00071[24] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [8] <= 1'h0;
      else \nr00071[24] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [9] <= 1'h0;
      else \nr00071[24] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [10] <= 1'h0;
      else \nr00071[24] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [11] <= 1'h0;
      else \nr00071[24] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [12] <= 1'h0;
      else \nr00071[24] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [13] <= 1'h0;
      else \nr00071[24] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [14] <= 1'h0;
      else \nr00071[24] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [15] <= 1'h0;
      else \nr00071[24] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [16] <= 1'h0;
      else \nr00071[24] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [17] <= 1'h0;
      else \nr00071[24] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [18] <= 1'h0;
      else \nr00071[24] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [19] <= 1'h0;
      else \nr00071[24] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [20] <= 1'h0;
      else \nr00071[24] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [21] <= 1'h0;
      else \nr00071[24] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [22] <= 1'h0;
      else \nr00071[24] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [23] <= 1'h0;
      else \nr00071[24] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [24] <= 1'h0;
      else \nr00071[24] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [25] <= 1'h0;
      else \nr00071[24] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [26] <= 1'h0;
      else \nr00071[24] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [27] <= 1'h0;
      else \nr00071[24] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [28] <= 1'h0;
      else \nr00071[24] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [29] <= 1'h0;
      else \nr00071[24] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [30] <= 1'h0;
      else \nr00071[24] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00024)
      if (!nw00400) \nr00071[24] [31] <= 1'h0;
      else \nr00071[24] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [0] <= 1'h0;
      else \nr00071[23] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [1] <= 1'h0;
      else \nr00071[23] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [2] <= 1'h0;
      else \nr00071[23] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [3] <= 1'h0;
      else \nr00071[23] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [4] <= 1'h0;
      else \nr00071[23] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [5] <= 1'h0;
      else \nr00071[23] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [6] <= 1'h0;
      else \nr00071[23] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [7] <= 1'h0;
      else \nr00071[23] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [8] <= 1'h0;
      else \nr00071[23] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [9] <= 1'h0;
      else \nr00071[23] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [10] <= 1'h0;
      else \nr00071[23] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [11] <= 1'h0;
      else \nr00071[23] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [12] <= 1'h0;
      else \nr00071[23] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [13] <= 1'h0;
      else \nr00071[23] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [14] <= 1'h0;
      else \nr00071[23] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [15] <= 1'h0;
      else \nr00071[23] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [16] <= 1'h0;
      else \nr00071[23] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [17] <= 1'h0;
      else \nr00071[23] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [18] <= 1'h0;
      else \nr00071[23] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [19] <= 1'h0;
      else \nr00071[23] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [20] <= 1'h0;
      else \nr00071[23] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [21] <= 1'h0;
      else \nr00071[23] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [22] <= 1'h0;
      else \nr00071[23] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [23] <= 1'h0;
      else \nr00071[23] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [24] <= 1'h0;
      else \nr00071[23] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [25] <= 1'h0;
      else \nr00071[23] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [26] <= 1'h0;
      else \nr00071[23] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [27] <= 1'h0;
      else \nr00071[23] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [28] <= 1'h0;
      else \nr00071[23] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [29] <= 1'h0;
      else \nr00071[23] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [30] <= 1'h0;
      else \nr00071[23] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00025)
      if (!nw00399) \nr00071[23] [31] <= 1'h0;
      else \nr00071[23] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [0] <= 1'h0;
      else \nr00071[22] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [1] <= 1'h0;
      else \nr00071[22] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [2] <= 1'h0;
      else \nr00071[22] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [3] <= 1'h0;
      else \nr00071[22] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [4] <= 1'h0;
      else \nr00071[22] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [5] <= 1'h0;
      else \nr00071[22] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [6] <= 1'h0;
      else \nr00071[22] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [7] <= 1'h0;
      else \nr00071[22] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [8] <= 1'h0;
      else \nr00071[22] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [9] <= 1'h0;
      else \nr00071[22] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [10] <= 1'h0;
      else \nr00071[22] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [11] <= 1'h0;
      else \nr00071[22] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [12] <= 1'h0;
      else \nr00071[22] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [13] <= 1'h0;
      else \nr00071[22] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [14] <= 1'h0;
      else \nr00071[22] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [15] <= 1'h0;
      else \nr00071[22] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [16] <= 1'h0;
      else \nr00071[22] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [17] <= 1'h0;
      else \nr00071[22] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [18] <= 1'h0;
      else \nr00071[22] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [19] <= 1'h0;
      else \nr00071[22] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [20] <= 1'h0;
      else \nr00071[22] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [21] <= 1'h0;
      else \nr00071[22] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [22] <= 1'h0;
      else \nr00071[22] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [23] <= 1'h0;
      else \nr00071[22] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [24] <= 1'h0;
      else \nr00071[22] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [25] <= 1'h0;
      else \nr00071[22] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [26] <= 1'h0;
      else \nr00071[22] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [27] <= 1'h0;
      else \nr00071[22] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [28] <= 1'h0;
      else \nr00071[22] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [29] <= 1'h0;
      else \nr00071[22] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [30] <= 1'h0;
      else \nr00071[22] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00026)
      if (!nw00398) \nr00071[22] [31] <= 1'h0;
      else \nr00071[22] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [0] <= 1'h0;
      else \nr00071[21] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [1] <= 1'h0;
      else \nr00071[21] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [2] <= 1'h0;
      else \nr00071[21] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [3] <= 1'h0;
      else \nr00071[21] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [4] <= 1'h0;
      else \nr00071[21] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [5] <= 1'h0;
      else \nr00071[21] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [6] <= 1'h0;
      else \nr00071[21] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [7] <= 1'h0;
      else \nr00071[21] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [8] <= 1'h0;
      else \nr00071[21] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [9] <= 1'h0;
      else \nr00071[21] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [10] <= 1'h0;
      else \nr00071[21] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [11] <= 1'h0;
      else \nr00071[21] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [12] <= 1'h0;
      else \nr00071[21] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [13] <= 1'h0;
      else \nr00071[21] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [14] <= 1'h0;
      else \nr00071[21] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [15] <= 1'h0;
      else \nr00071[21] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [16] <= 1'h0;
      else \nr00071[21] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [17] <= 1'h0;
      else \nr00071[21] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [18] <= 1'h0;
      else \nr00071[21] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [19] <= 1'h0;
      else \nr00071[21] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [20] <= 1'h0;
      else \nr00071[21] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [21] <= 1'h0;
      else \nr00071[21] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [22] <= 1'h0;
      else \nr00071[21] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [23] <= 1'h0;
      else \nr00071[21] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [24] <= 1'h0;
      else \nr00071[21] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [25] <= 1'h0;
      else \nr00071[21] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [26] <= 1'h0;
      else \nr00071[21] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [27] <= 1'h0;
      else \nr00071[21] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [28] <= 1'h0;
      else \nr00071[21] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [29] <= 1'h0;
      else \nr00071[21] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [30] <= 1'h0;
      else \nr00071[21] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00027)
      if (!nw00397) \nr00071[21] [31] <= 1'h0;
      else \nr00071[21] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [0] <= 1'h0;
      else \nr00071[20] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [1] <= 1'h0;
      else \nr00071[20] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [2] <= 1'h0;
      else \nr00071[20] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [3] <= 1'h0;
      else \nr00071[20] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [4] <= 1'h0;
      else \nr00071[20] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [5] <= 1'h0;
      else \nr00071[20] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [6] <= 1'h0;
      else \nr00071[20] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [7] <= 1'h0;
      else \nr00071[20] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [8] <= 1'h0;
      else \nr00071[20] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [9] <= 1'h0;
      else \nr00071[20] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [10] <= 1'h0;
      else \nr00071[20] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [11] <= 1'h0;
      else \nr00071[20] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [12] <= 1'h0;
      else \nr00071[20] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [13] <= 1'h0;
      else \nr00071[20] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [14] <= 1'h0;
      else \nr00071[20] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [15] <= 1'h0;
      else \nr00071[20] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [16] <= 1'h0;
      else \nr00071[20] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [17] <= 1'h0;
      else \nr00071[20] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [18] <= 1'h0;
      else \nr00071[20] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [19] <= 1'h0;
      else \nr00071[20] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [20] <= 1'h0;
      else \nr00071[20] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [21] <= 1'h0;
      else \nr00071[20] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [22] <= 1'h0;
      else \nr00071[20] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [23] <= 1'h0;
      else \nr00071[20] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [24] <= 1'h0;
      else \nr00071[20] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [25] <= 1'h0;
      else \nr00071[20] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [26] <= 1'h0;
      else \nr00071[20] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [27] <= 1'h0;
      else \nr00071[20] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [28] <= 1'h0;
      else \nr00071[20] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [29] <= 1'h0;
      else \nr00071[20] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [30] <= 1'h0;
      else \nr00071[20] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00028)
      if (!nw00396) \nr00071[20] [31] <= 1'h0;
      else \nr00071[20] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [0] <= 1'h0;
      else \nr00071[19] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [1] <= 1'h0;
      else \nr00071[19] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [2] <= 1'h0;
      else \nr00071[19] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [3] <= 1'h0;
      else \nr00071[19] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [4] <= 1'h0;
      else \nr00071[19] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [5] <= 1'h0;
      else \nr00071[19] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [6] <= 1'h0;
      else \nr00071[19] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [7] <= 1'h0;
      else \nr00071[19] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [8] <= 1'h0;
      else \nr00071[19] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [9] <= 1'h0;
      else \nr00071[19] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [10] <= 1'h0;
      else \nr00071[19] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [11] <= 1'h0;
      else \nr00071[19] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [12] <= 1'h0;
      else \nr00071[19] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [13] <= 1'h0;
      else \nr00071[19] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [14] <= 1'h0;
      else \nr00071[19] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [15] <= 1'h0;
      else \nr00071[19] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [16] <= 1'h0;
      else \nr00071[19] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [17] <= 1'h0;
      else \nr00071[19] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [18] <= 1'h0;
      else \nr00071[19] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [19] <= 1'h0;
      else \nr00071[19] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [20] <= 1'h0;
      else \nr00071[19] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [21] <= 1'h0;
      else \nr00071[19] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [22] <= 1'h0;
      else \nr00071[19] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [23] <= 1'h0;
      else \nr00071[19] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [24] <= 1'h0;
      else \nr00071[19] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [25] <= 1'h0;
      else \nr00071[19] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [26] <= 1'h0;
      else \nr00071[19] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [27] <= 1'h0;
      else \nr00071[19] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [28] <= 1'h0;
      else \nr00071[19] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [29] <= 1'h0;
      else \nr00071[19] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [30] <= 1'h0;
      else \nr00071[19] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00030)
      if (!nw00394) \nr00071[19] [31] <= 1'h0;
      else \nr00071[19] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [0] <= 1'h0;
      else \nr00071[18] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [1] <= 1'h0;
      else \nr00071[18] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [2] <= 1'h0;
      else \nr00071[18] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [3] <= 1'h0;
      else \nr00071[18] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [4] <= 1'h0;
      else \nr00071[18] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [5] <= 1'h0;
      else \nr00071[18] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [6] <= 1'h0;
      else \nr00071[18] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [7] <= 1'h0;
      else \nr00071[18] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [8] <= 1'h0;
      else \nr00071[18] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [9] <= 1'h0;
      else \nr00071[18] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [10] <= 1'h0;
      else \nr00071[18] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [11] <= 1'h0;
      else \nr00071[18] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [12] <= 1'h0;
      else \nr00071[18] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [13] <= 1'h0;
      else \nr00071[18] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [14] <= 1'h0;
      else \nr00071[18] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [15] <= 1'h0;
      else \nr00071[18] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [16] <= 1'h0;
      else \nr00071[18] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [17] <= 1'h0;
      else \nr00071[18] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [18] <= 1'h0;
      else \nr00071[18] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [19] <= 1'h0;
      else \nr00071[18] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [20] <= 1'h0;
      else \nr00071[18] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [21] <= 1'h0;
      else \nr00071[18] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [22] <= 1'h0;
      else \nr00071[18] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [23] <= 1'h0;
      else \nr00071[18] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [24] <= 1'h0;
      else \nr00071[18] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [25] <= 1'h0;
      else \nr00071[18] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [26] <= 1'h0;
      else \nr00071[18] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [27] <= 1'h0;
      else \nr00071[18] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [28] <= 1'h0;
      else \nr00071[18] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [29] <= 1'h0;
      else \nr00071[18] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [30] <= 1'h0;
      else \nr00071[18] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00031)
      if (!nw00393) \nr00071[18] [31] <= 1'h0;
      else \nr00071[18] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [0] <= 1'h0;
      else \nr00071[17] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [1] <= 1'h0;
      else \nr00071[17] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [2] <= 1'h0;
      else \nr00071[17] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [3] <= 1'h0;
      else \nr00071[17] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [4] <= 1'h0;
      else \nr00071[17] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [5] <= 1'h0;
      else \nr00071[17] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [6] <= 1'h0;
      else \nr00071[17] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [7] <= 1'h0;
      else \nr00071[17] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [8] <= 1'h0;
      else \nr00071[17] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [9] <= 1'h0;
      else \nr00071[17] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [10] <= 1'h0;
      else \nr00071[17] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [11] <= 1'h0;
      else \nr00071[17] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [12] <= 1'h0;
      else \nr00071[17] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [13] <= 1'h0;
      else \nr00071[17] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [14] <= 1'h0;
      else \nr00071[17] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [15] <= 1'h0;
      else \nr00071[17] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [16] <= 1'h0;
      else \nr00071[17] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [17] <= 1'h0;
      else \nr00071[17] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [18] <= 1'h0;
      else \nr00071[17] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [19] <= 1'h0;
      else \nr00071[17] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [20] <= 1'h0;
      else \nr00071[17] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [21] <= 1'h0;
      else \nr00071[17] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [22] <= 1'h0;
      else \nr00071[17] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [23] <= 1'h0;
      else \nr00071[17] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [24] <= 1'h0;
      else \nr00071[17] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [25] <= 1'h0;
      else \nr00071[17] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [26] <= 1'h0;
      else \nr00071[17] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [27] <= 1'h0;
      else \nr00071[17] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [28] <= 1'h0;
      else \nr00071[17] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [29] <= 1'h0;
      else \nr00071[17] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [30] <= 1'h0;
      else \nr00071[17] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00032)
      if (!nw00392) \nr00071[17] [31] <= 1'h0;
      else \nr00071[17] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [0] <= 1'h0;
      else \nr00071[16] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [1] <= 1'h0;
      else \nr00071[16] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [2] <= 1'h0;
      else \nr00071[16] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [3] <= 1'h0;
      else \nr00071[16] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [4] <= 1'h0;
      else \nr00071[16] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [5] <= 1'h0;
      else \nr00071[16] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [6] <= 1'h0;
      else \nr00071[16] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [7] <= 1'h0;
      else \nr00071[16] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [8] <= 1'h0;
      else \nr00071[16] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [9] <= 1'h0;
      else \nr00071[16] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [10] <= 1'h0;
      else \nr00071[16] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [11] <= 1'h0;
      else \nr00071[16] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [12] <= 1'h0;
      else \nr00071[16] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [13] <= 1'h0;
      else \nr00071[16] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [14] <= 1'h0;
      else \nr00071[16] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [15] <= 1'h0;
      else \nr00071[16] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [16] <= 1'h0;
      else \nr00071[16] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [17] <= 1'h0;
      else \nr00071[16] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [18] <= 1'h0;
      else \nr00071[16] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [19] <= 1'h0;
      else \nr00071[16] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [20] <= 1'h0;
      else \nr00071[16] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [21] <= 1'h0;
      else \nr00071[16] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [22] <= 1'h0;
      else \nr00071[16] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [23] <= 1'h0;
      else \nr00071[16] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [24] <= 1'h0;
      else \nr00071[16] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [25] <= 1'h0;
      else \nr00071[16] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [26] <= 1'h0;
      else \nr00071[16] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [27] <= 1'h0;
      else \nr00071[16] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [28] <= 1'h0;
      else \nr00071[16] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [29] <= 1'h0;
      else \nr00071[16] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [30] <= 1'h0;
      else \nr00071[16] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00033)
      if (!nw00391) \nr00071[16] [31] <= 1'h0;
      else \nr00071[16] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [0] <= 1'h0;
      else \nr00071[15] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [1] <= 1'h0;
      else \nr00071[15] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [2] <= 1'h0;
      else \nr00071[15] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [3] <= 1'h0;
      else \nr00071[15] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [4] <= 1'h0;
      else \nr00071[15] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [5] <= 1'h0;
      else \nr00071[15] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [6] <= 1'h0;
      else \nr00071[15] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [7] <= 1'h0;
      else \nr00071[15] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [8] <= 1'h0;
      else \nr00071[15] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [9] <= 1'h0;
      else \nr00071[15] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [10] <= 1'h0;
      else \nr00071[15] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [11] <= 1'h0;
      else \nr00071[15] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [12] <= 1'h0;
      else \nr00071[15] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [13] <= 1'h0;
      else \nr00071[15] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [14] <= 1'h0;
      else \nr00071[15] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [15] <= 1'h0;
      else \nr00071[15] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [16] <= 1'h0;
      else \nr00071[15] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [17] <= 1'h0;
      else \nr00071[15] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [18] <= 1'h0;
      else \nr00071[15] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [19] <= 1'h0;
      else \nr00071[15] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [20] <= 1'h0;
      else \nr00071[15] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [21] <= 1'h0;
      else \nr00071[15] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [22] <= 1'h0;
      else \nr00071[15] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [23] <= 1'h0;
      else \nr00071[15] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [24] <= 1'h0;
      else \nr00071[15] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [25] <= 1'h0;
      else \nr00071[15] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [26] <= 1'h0;
      else \nr00071[15] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [27] <= 1'h0;
      else \nr00071[15] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [28] <= 1'h0;
      else \nr00071[15] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [29] <= 1'h0;
      else \nr00071[15] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [30] <= 1'h0;
      else \nr00071[15] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00034)
      if (!nw00390) \nr00071[15] [31] <= 1'h0;
      else \nr00071[15] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [0] <= 1'h0;
      else \nr00071[14] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [1] <= 1'h0;
      else \nr00071[14] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [2] <= 1'h0;
      else \nr00071[14] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [3] <= 1'h0;
      else \nr00071[14] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [4] <= 1'h0;
      else \nr00071[14] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [5] <= 1'h0;
      else \nr00071[14] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [6] <= 1'h0;
      else \nr00071[14] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [7] <= 1'h0;
      else \nr00071[14] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [8] <= 1'h0;
      else \nr00071[14] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [9] <= 1'h0;
      else \nr00071[14] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [10] <= 1'h0;
      else \nr00071[14] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [11] <= 1'h0;
      else \nr00071[14] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [12] <= 1'h0;
      else \nr00071[14] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [13] <= 1'h0;
      else \nr00071[14] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [14] <= 1'h0;
      else \nr00071[14] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [15] <= 1'h0;
      else \nr00071[14] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [16] <= 1'h0;
      else \nr00071[14] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [17] <= 1'h0;
      else \nr00071[14] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [18] <= 1'h0;
      else \nr00071[14] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [19] <= 1'h0;
      else \nr00071[14] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [20] <= 1'h0;
      else \nr00071[14] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [21] <= 1'h0;
      else \nr00071[14] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [22] <= 1'h0;
      else \nr00071[14] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [23] <= 1'h0;
      else \nr00071[14] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [24] <= 1'h0;
      else \nr00071[14] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [25] <= 1'h0;
      else \nr00071[14] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [26] <= 1'h0;
      else \nr00071[14] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [27] <= 1'h0;
      else \nr00071[14] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [28] <= 1'h0;
      else \nr00071[14] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [29] <= 1'h0;
      else \nr00071[14] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [30] <= 1'h0;
      else \nr00071[14] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00035)
      if (!nw00389) \nr00071[14] [31] <= 1'h0;
      else \nr00071[14] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [0] <= 1'h0;
      else \nr00071[13] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [1] <= 1'h0;
      else \nr00071[13] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [2] <= 1'h0;
      else \nr00071[13] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [3] <= 1'h0;
      else \nr00071[13] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [4] <= 1'h0;
      else \nr00071[13] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [5] <= 1'h0;
      else \nr00071[13] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [6] <= 1'h0;
      else \nr00071[13] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [7] <= 1'h0;
      else \nr00071[13] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [8] <= 1'h0;
      else \nr00071[13] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [9] <= 1'h0;
      else \nr00071[13] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [10] <= 1'h0;
      else \nr00071[13] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [11] <= 1'h0;
      else \nr00071[13] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [12] <= 1'h0;
      else \nr00071[13] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [13] <= 1'h0;
      else \nr00071[13] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [14] <= 1'h0;
      else \nr00071[13] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [15] <= 1'h0;
      else \nr00071[13] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [16] <= 1'h0;
      else \nr00071[13] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [17] <= 1'h0;
      else \nr00071[13] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [18] <= 1'h0;
      else \nr00071[13] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [19] <= 1'h0;
      else \nr00071[13] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [20] <= 1'h0;
      else \nr00071[13] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [21] <= 1'h0;
      else \nr00071[13] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [22] <= 1'h0;
      else \nr00071[13] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [23] <= 1'h0;
      else \nr00071[13] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [24] <= 1'h0;
      else \nr00071[13] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [25] <= 1'h0;
      else \nr00071[13] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [26] <= 1'h0;
      else \nr00071[13] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [27] <= 1'h0;
      else \nr00071[13] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [28] <= 1'h0;
      else \nr00071[13] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [29] <= 1'h0;
      else \nr00071[13] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [30] <= 1'h0;
      else \nr00071[13] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00036)
      if (!nw00388) \nr00071[13] [31] <= 1'h0;
      else \nr00071[13] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [0] <= 1'h0;
      else \nr00071[12] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [1] <= 1'h0;
      else \nr00071[12] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [2] <= 1'h0;
      else \nr00071[12] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [3] <= 1'h0;
      else \nr00071[12] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [4] <= 1'h0;
      else \nr00071[12] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [5] <= 1'h0;
      else \nr00071[12] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [6] <= 1'h0;
      else \nr00071[12] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [7] <= 1'h0;
      else \nr00071[12] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [8] <= 1'h0;
      else \nr00071[12] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [9] <= 1'h0;
      else \nr00071[12] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [10] <= 1'h0;
      else \nr00071[12] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [11] <= 1'h0;
      else \nr00071[12] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [12] <= 1'h0;
      else \nr00071[12] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [13] <= 1'h0;
      else \nr00071[12] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [14] <= 1'h0;
      else \nr00071[12] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [15] <= 1'h0;
      else \nr00071[12] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [16] <= 1'h0;
      else \nr00071[12] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [17] <= 1'h0;
      else \nr00071[12] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [18] <= 1'h0;
      else \nr00071[12] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [19] <= 1'h0;
      else \nr00071[12] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [20] <= 1'h0;
      else \nr00071[12] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [21] <= 1'h0;
      else \nr00071[12] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [22] <= 1'h0;
      else \nr00071[12] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [23] <= 1'h0;
      else \nr00071[12] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [24] <= 1'h0;
      else \nr00071[12] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [25] <= 1'h0;
      else \nr00071[12] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [26] <= 1'h0;
      else \nr00071[12] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [27] <= 1'h0;
      else \nr00071[12] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [28] <= 1'h0;
      else \nr00071[12] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [29] <= 1'h0;
      else \nr00071[12] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [30] <= 1'h0;
      else \nr00071[12] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00037)
      if (!nw00387) \nr00071[12] [31] <= 1'h0;
      else \nr00071[12] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [0] <= 1'h0;
      else \nr00071[11] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [1] <= 1'h0;
      else \nr00071[11] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [2] <= 1'h0;
      else \nr00071[11] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [3] <= 1'h0;
      else \nr00071[11] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [4] <= 1'h0;
      else \nr00071[11] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [5] <= 1'h0;
      else \nr00071[11] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [6] <= 1'h0;
      else \nr00071[11] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [7] <= 1'h0;
      else \nr00071[11] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [8] <= 1'h0;
      else \nr00071[11] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [9] <= 1'h0;
      else \nr00071[11] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [10] <= 1'h0;
      else \nr00071[11] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [11] <= 1'h0;
      else \nr00071[11] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [12] <= 1'h0;
      else \nr00071[11] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [13] <= 1'h0;
      else \nr00071[11] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [14] <= 1'h0;
      else \nr00071[11] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [15] <= 1'h0;
      else \nr00071[11] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [16] <= 1'h0;
      else \nr00071[11] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [17] <= 1'h0;
      else \nr00071[11] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [18] <= 1'h0;
      else \nr00071[11] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [19] <= 1'h0;
      else \nr00071[11] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [20] <= 1'h0;
      else \nr00071[11] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [21] <= 1'h0;
      else \nr00071[11] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [22] <= 1'h0;
      else \nr00071[11] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [23] <= 1'h0;
      else \nr00071[11] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [24] <= 1'h0;
      else \nr00071[11] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [25] <= 1'h0;
      else \nr00071[11] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [26] <= 1'h0;
      else \nr00071[11] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [27] <= 1'h0;
      else \nr00071[11] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [28] <= 1'h0;
      else \nr00071[11] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [29] <= 1'h0;
      else \nr00071[11] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [30] <= 1'h0;
      else \nr00071[11] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00038)
      if (!nw00386) \nr00071[11] [31] <= 1'h0;
      else \nr00071[11] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [0] <= 1'h0;
    else \nr00071[0] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [1] <= 1'h0;
    else \nr00071[0] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [2] <= 1'h0;
    else \nr00071[0] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [3] <= 1'h0;
    else \nr00071[0] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [4] <= 1'h0;
    else \nr00071[0] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [5] <= 1'h0;
    else \nr00071[0] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [6] <= 1'h0;
    else \nr00071[0] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [7] <= 1'h0;
    else \nr00071[0] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [8] <= 1'h0;
    else \nr00071[0] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [9] <= 1'h0;
    else \nr00071[0] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [10] <= 1'h0;
    else \nr00071[0] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [11] <= 1'h0;
    else \nr00071[0] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [12] <= 1'h0;
    else \nr00071[0] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [13] <= 1'h0;
    else \nr00071[0] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [14] <= 1'h0;
    else \nr00071[0] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [15] <= 1'h0;
    else \nr00071[0] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [16] <= 1'h0;
    else \nr00071[0] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [17] <= 1'h0;
    else \nr00071[0] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [18] <= 1'h0;
    else \nr00071[0] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [19] <= 1'h0;
    else \nr00071[0] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [20] <= 1'h0;
    else \nr00071[0] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [21] <= 1'h0;
    else \nr00071[0] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [22] <= 1'h0;
    else \nr00071[0] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [23] <= 1'h0;
    else \nr00071[0] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [24] <= 1'h0;
    else \nr00071[0] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [25] <= 1'h0;
    else \nr00071[0] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [26] <= 1'h0;
    else \nr00071[0] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [27] <= 1'h0;
    else \nr00071[0] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [28] <= 1'h0;
    else \nr00071[0] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [29] <= 1'h0;
    else \nr00071[0] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [30] <= 1'h0;
    else \nr00071[0] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (!nw00384) \nr00071[0] [31] <= 1'h0;
    else \nr00071[0] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [0] <= 1'h0;
      else \nr00071[9] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [1] <= 1'h0;
      else \nr00071[9] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [2] <= 1'h0;
      else \nr00071[9] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [3] <= 1'h0;
      else \nr00071[9] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [4] <= 1'h0;
      else \nr00071[9] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [5] <= 1'h0;
      else \nr00071[9] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [6] <= 1'h0;
      else \nr00071[9] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [7] <= 1'h0;
      else \nr00071[9] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [8] <= 1'h0;
      else \nr00071[9] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [9] <= 1'h0;
      else \nr00071[9] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [10] <= 1'h0;
      else \nr00071[9] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [11] <= 1'h0;
      else \nr00071[9] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [12] <= 1'h0;
      else \nr00071[9] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [13] <= 1'h0;
      else \nr00071[9] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [14] <= 1'h0;
      else \nr00071[9] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [15] <= 1'h0;
      else \nr00071[9] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [16] <= 1'h0;
      else \nr00071[9] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [17] <= 1'h0;
      else \nr00071[9] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [18] <= 1'h0;
      else \nr00071[9] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [19] <= 1'h0;
      else \nr00071[9] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [20] <= 1'h0;
      else \nr00071[9] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [21] <= 1'h0;
      else \nr00071[9] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [22] <= 1'h0;
      else \nr00071[9] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [23] <= 1'h0;
      else \nr00071[9] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [24] <= 1'h0;
      else \nr00071[9] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [25] <= 1'h0;
      else \nr00071[9] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [26] <= 1'h0;
      else \nr00071[9] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [27] <= 1'h0;
      else \nr00071[9] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [28] <= 1'h0;
      else \nr00071[9] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [29] <= 1'h0;
      else \nr00071[9] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [30] <= 1'h0;
      else \nr00071[9] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00009)
      if (!nw00415) \nr00071[9] [31] <= 1'h0;
      else \nr00071[9] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [0] <= 1'h0;
      else \nr00071[8] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [1] <= 1'h0;
      else \nr00071[8] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [2] <= 1'h0;
      else \nr00071[8] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [3] <= 1'h0;
      else \nr00071[8] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [4] <= 1'h0;
      else \nr00071[8] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [5] <= 1'h0;
      else \nr00071[8] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [6] <= 1'h0;
      else \nr00071[8] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [7] <= 1'h0;
      else \nr00071[8] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [8] <= 1'h0;
      else \nr00071[8] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [9] <= 1'h0;
      else \nr00071[8] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [10] <= 1'h0;
      else \nr00071[8] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [11] <= 1'h0;
      else \nr00071[8] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [12] <= 1'h0;
      else \nr00071[8] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [13] <= 1'h0;
      else \nr00071[8] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [14] <= 1'h0;
      else \nr00071[8] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [15] <= 1'h0;
      else \nr00071[8] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [16] <= 1'h0;
      else \nr00071[8] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [17] <= 1'h0;
      else \nr00071[8] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [18] <= 1'h0;
      else \nr00071[8] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [19] <= 1'h0;
      else \nr00071[8] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [20] <= 1'h0;
      else \nr00071[8] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [21] <= 1'h0;
      else \nr00071[8] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [22] <= 1'h0;
      else \nr00071[8] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [23] <= 1'h0;
      else \nr00071[8] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [24] <= 1'h0;
      else \nr00071[8] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [25] <= 1'h0;
      else \nr00071[8] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [26] <= 1'h0;
      else \nr00071[8] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [27] <= 1'h0;
      else \nr00071[8] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [28] <= 1'h0;
      else \nr00071[8] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [29] <= 1'h0;
      else \nr00071[8] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [30] <= 1'h0;
      else \nr00071[8] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00010)
      if (!nw00414) \nr00071[8] [31] <= 1'h0;
      else \nr00071[8] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [0] <= 1'h0;
      else \nr00071[7] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [1] <= 1'h0;
      else \nr00071[7] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [2] <= 1'h0;
      else \nr00071[7] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [3] <= 1'h0;
      else \nr00071[7] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [4] <= 1'h0;
      else \nr00071[7] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [5] <= 1'h0;
      else \nr00071[7] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [6] <= 1'h0;
      else \nr00071[7] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [7] <= 1'h0;
      else \nr00071[7] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [8] <= 1'h0;
      else \nr00071[7] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [9] <= 1'h0;
      else \nr00071[7] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [10] <= 1'h0;
      else \nr00071[7] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [11] <= 1'h0;
      else \nr00071[7] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [12] <= 1'h0;
      else \nr00071[7] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [13] <= 1'h0;
      else \nr00071[7] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [14] <= 1'h0;
      else \nr00071[7] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [15] <= 1'h0;
      else \nr00071[7] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [16] <= 1'h0;
      else \nr00071[7] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [17] <= 1'h0;
      else \nr00071[7] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [18] <= 1'h0;
      else \nr00071[7] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [19] <= 1'h0;
      else \nr00071[7] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [20] <= 1'h0;
      else \nr00071[7] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [21] <= 1'h0;
      else \nr00071[7] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [22] <= 1'h0;
      else \nr00071[7] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [23] <= 1'h0;
      else \nr00071[7] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [24] <= 1'h0;
      else \nr00071[7] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [25] <= 1'h0;
      else \nr00071[7] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [26] <= 1'h0;
      else \nr00071[7] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [27] <= 1'h0;
      else \nr00071[7] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [28] <= 1'h0;
      else \nr00071[7] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [29] <= 1'h0;
      else \nr00071[7] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [30] <= 1'h0;
      else \nr00071[7] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00011)
      if (!nw00413) \nr00071[7] [31] <= 1'h0;
      else \nr00071[7] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [0] <= 1'h0;
      else \nr00071[6] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [1] <= 1'h0;
      else \nr00071[6] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [2] <= 1'h0;
      else \nr00071[6] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [3] <= 1'h0;
      else \nr00071[6] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [4] <= 1'h0;
      else \nr00071[6] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [5] <= 1'h0;
      else \nr00071[6] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [6] <= 1'h0;
      else \nr00071[6] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [7] <= 1'h0;
      else \nr00071[6] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [8] <= 1'h0;
      else \nr00071[6] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [9] <= 1'h0;
      else \nr00071[6] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [10] <= 1'h0;
      else \nr00071[6] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [11] <= 1'h0;
      else \nr00071[6] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [12] <= 1'h0;
      else \nr00071[6] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [13] <= 1'h0;
      else \nr00071[6] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [14] <= 1'h0;
      else \nr00071[6] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [15] <= 1'h0;
      else \nr00071[6] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [16] <= 1'h0;
      else \nr00071[6] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [17] <= 1'h0;
      else \nr00071[6] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [18] <= 1'h0;
      else \nr00071[6] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [19] <= 1'h0;
      else \nr00071[6] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [20] <= 1'h0;
      else \nr00071[6] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [21] <= 1'h0;
      else \nr00071[6] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [22] <= 1'h0;
      else \nr00071[6] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [23] <= 1'h0;
      else \nr00071[6] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [24] <= 1'h0;
      else \nr00071[6] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [25] <= 1'h0;
      else \nr00071[6] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [26] <= 1'h0;
      else \nr00071[6] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [27] <= 1'h0;
      else \nr00071[6] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [28] <= 1'h0;
      else \nr00071[6] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [29] <= 1'h0;
      else \nr00071[6] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [30] <= 1'h0;
      else \nr00071[6] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00012)
      if (!nw00412) \nr00071[6] [31] <= 1'h0;
      else \nr00071[6] [31] <= nw00089;
  always @(posedge clock_10_i)
    nr00000[0] <= nw00055;
  always @(posedge clock_10_i)
    nr00000[1] <= nw00056;
  always @(posedge clock_10_i)
    nr00000[2] <= nw00057;
  always @(posedge clock_10_i)
    nr00000[3] <= nw00058;
  always @(posedge clock_10_i)
    nr00000[4] <= nw00059;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [0] <= 1'h0;
      else \nr00071[31] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [1] <= 1'h0;
      else \nr00071[31] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [2] <= 1'h0;
      else \nr00071[31] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [3] <= 1'h0;
      else \nr00071[31] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [4] <= 1'h0;
      else \nr00071[31] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [5] <= 1'h0;
      else \nr00071[31] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [6] <= 1'h0;
      else \nr00071[31] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [7] <= 1'h0;
      else \nr00071[31] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [8] <= 1'h0;
      else \nr00071[31] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [9] <= 1'h0;
      else \nr00071[31] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [10] <= 1'h0;
      else \nr00071[31] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [11] <= 1'h0;
      else \nr00071[31] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [12] <= 1'h0;
      else \nr00071[31] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [13] <= 1'h0;
      else \nr00071[31] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [14] <= 1'h0;
      else \nr00071[31] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [15] <= 1'h0;
      else \nr00071[31] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [16] <= 1'h0;
      else \nr00071[31] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [17] <= 1'h0;
      else \nr00071[31] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [18] <= 1'h0;
      else \nr00071[31] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [19] <= 1'h0;
      else \nr00071[31] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [20] <= 1'h0;
      else \nr00071[31] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [21] <= 1'h0;
      else \nr00071[31] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [22] <= 1'h0;
      else \nr00071[31] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [23] <= 1'h0;
      else \nr00071[31] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [24] <= 1'h0;
      else \nr00071[31] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [25] <= 1'h0;
      else \nr00071[31] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [26] <= 1'h0;
      else \nr00071[31] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [27] <= 1'h0;
      else \nr00071[31] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [28] <= 1'h0;
      else \nr00071[31] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [29] <= 1'h0;
      else \nr00071[31] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [30] <= 1'h0;
      else \nr00071[31] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00016)
      if (!nw00408) \nr00071[31] [31] <= 1'h0;
      else \nr00071[31] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [0] <= 1'h0;
      else \nr00071[5] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [1] <= 1'h0;
      else \nr00071[5] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [2] <= 1'h0;
      else \nr00071[5] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [3] <= 1'h0;
      else \nr00071[5] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [4] <= 1'h0;
      else \nr00071[5] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [5] <= 1'h0;
      else \nr00071[5] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [6] <= 1'h0;
      else \nr00071[5] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [7] <= 1'h0;
      else \nr00071[5] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [8] <= 1'h0;
      else \nr00071[5] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [9] <= 1'h0;
      else \nr00071[5] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [10] <= 1'h0;
      else \nr00071[5] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [11] <= 1'h0;
      else \nr00071[5] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [12] <= 1'h0;
      else \nr00071[5] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [13] <= 1'h0;
      else \nr00071[5] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [14] <= 1'h0;
      else \nr00071[5] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [15] <= 1'h0;
      else \nr00071[5] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [16] <= 1'h0;
      else \nr00071[5] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [17] <= 1'h0;
      else \nr00071[5] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [18] <= 1'h0;
      else \nr00071[5] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [19] <= 1'h0;
      else \nr00071[5] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [20] <= 1'h0;
      else \nr00071[5] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [21] <= 1'h0;
      else \nr00071[5] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [22] <= 1'h0;
      else \nr00071[5] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [23] <= 1'h0;
      else \nr00071[5] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [24] <= 1'h0;
      else \nr00071[5] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [25] <= 1'h0;
      else \nr00071[5] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [26] <= 1'h0;
      else \nr00071[5] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [27] <= 1'h0;
      else \nr00071[5] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [28] <= 1'h0;
      else \nr00071[5] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [29] <= 1'h0;
      else \nr00071[5] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [30] <= 1'h0;
      else \nr00071[5] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00013)
      if (!nw00411) \nr00071[5] [31] <= 1'h0;
      else \nr00071[5] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [0] <= 1'h0;
      else \nr00071[4] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [1] <= 1'h0;
      else \nr00071[4] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [2] <= 1'h0;
      else \nr00071[4] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [3] <= 1'h0;
      else \nr00071[4] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [4] <= 1'h0;
      else \nr00071[4] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [5] <= 1'h0;
      else \nr00071[4] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [6] <= 1'h0;
      else \nr00071[4] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [7] <= 1'h0;
      else \nr00071[4] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [8] <= 1'h0;
      else \nr00071[4] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [9] <= 1'h0;
      else \nr00071[4] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [10] <= 1'h0;
      else \nr00071[4] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [11] <= 1'h0;
      else \nr00071[4] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [12] <= 1'h0;
      else \nr00071[4] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [13] <= 1'h0;
      else \nr00071[4] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [14] <= 1'h0;
      else \nr00071[4] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [15] <= 1'h0;
      else \nr00071[4] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [16] <= 1'h0;
      else \nr00071[4] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [17] <= 1'h0;
      else \nr00071[4] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [18] <= 1'h0;
      else \nr00071[4] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [19] <= 1'h0;
      else \nr00071[4] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [20] <= 1'h0;
      else \nr00071[4] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [21] <= 1'h0;
      else \nr00071[4] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [22] <= 1'h0;
      else \nr00071[4] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [23] <= 1'h0;
      else \nr00071[4] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [24] <= 1'h0;
      else \nr00071[4] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [25] <= 1'h0;
      else \nr00071[4] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [26] <= 1'h0;
      else \nr00071[4] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [27] <= 1'h0;
      else \nr00071[4] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [28] <= 1'h0;
      else \nr00071[4] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [29] <= 1'h0;
      else \nr00071[4] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [30] <= 1'h0;
      else \nr00071[4] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00014)
      if (!nw00410) \nr00071[4] [31] <= 1'h0;
      else \nr00071[4] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [0] <= 1'h0;
      else \nr00071[3] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [1] <= 1'h0;
      else \nr00071[3] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [2] <= 1'h0;
      else \nr00071[3] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [3] <= 1'h0;
      else \nr00071[3] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [4] <= 1'h0;
      else \nr00071[3] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [5] <= 1'h0;
      else \nr00071[3] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [6] <= 1'h0;
      else \nr00071[3] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [7] <= 1'h0;
      else \nr00071[3] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [8] <= 1'h0;
      else \nr00071[3] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [9] <= 1'h0;
      else \nr00071[3] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [10] <= 1'h0;
      else \nr00071[3] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [11] <= 1'h0;
      else \nr00071[3] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [12] <= 1'h0;
      else \nr00071[3] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [13] <= 1'h0;
      else \nr00071[3] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [14] <= 1'h0;
      else \nr00071[3] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [15] <= 1'h0;
      else \nr00071[3] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [16] <= 1'h0;
      else \nr00071[3] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [17] <= 1'h0;
      else \nr00071[3] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [18] <= 1'h0;
      else \nr00071[3] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [19] <= 1'h0;
      else \nr00071[3] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [20] <= 1'h0;
      else \nr00071[3] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [21] <= 1'h0;
      else \nr00071[3] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [22] <= 1'h0;
      else \nr00071[3] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [23] <= 1'h0;
      else \nr00071[3] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [24] <= 1'h0;
      else \nr00071[3] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [25] <= 1'h0;
      else \nr00071[3] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [26] <= 1'h0;
      else \nr00071[3] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [27] <= 1'h0;
      else \nr00071[3] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [28] <= 1'h0;
      else \nr00071[3] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [29] <= 1'h0;
      else \nr00071[3] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [30] <= 1'h0;
      else \nr00071[3] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00015)
      if (!nw00409) \nr00071[3] [31] <= 1'h0;
      else \nr00071[3] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [0] <= 1'h0;
      else \nr00071[2] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [1] <= 1'h0;
      else \nr00071[2] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [2] <= 1'h0;
      else \nr00071[2] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [3] <= 1'h0;
      else \nr00071[2] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [4] <= 1'h0;
      else \nr00071[2] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [5] <= 1'h0;
      else \nr00071[2] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [6] <= 1'h0;
      else \nr00071[2] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [7] <= 1'h0;
      else \nr00071[2] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [8] <= 1'h0;
      else \nr00071[2] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [9] <= 1'h0;
      else \nr00071[2] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [10] <= 1'h0;
      else \nr00071[2] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [11] <= 1'h0;
      else \nr00071[2] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [12] <= 1'h0;
      else \nr00071[2] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [13] <= 1'h0;
      else \nr00071[2] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [14] <= 1'h0;
      else \nr00071[2] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [15] <= 1'h0;
      else \nr00071[2] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [16] <= 1'h0;
      else \nr00071[2] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [17] <= 1'h0;
      else \nr00071[2] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [18] <= 1'h0;
      else \nr00071[2] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [19] <= 1'h0;
      else \nr00071[2] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [20] <= 1'h0;
      else \nr00071[2] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [21] <= 1'h0;
      else \nr00071[2] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [22] <= 1'h0;
      else \nr00071[2] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [23] <= 1'h0;
      else \nr00071[2] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [24] <= 1'h0;
      else \nr00071[2] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [25] <= 1'h0;
      else \nr00071[2] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [26] <= 1'h0;
      else \nr00071[2] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [27] <= 1'h0;
      else \nr00071[2] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [28] <= 1'h0;
      else \nr00071[2] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [29] <= 1'h0;
      else \nr00071[2] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [30] <= 1'h0;
      else \nr00071[2] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00018)
      if (!nw00406) \nr00071[2] [31] <= 1'h0;
      else \nr00071[2] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [0] <= 1'h0;
      else \nr00071[1] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [1] <= 1'h0;
      else \nr00071[1] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [2] <= 1'h0;
      else \nr00071[1] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [3] <= 1'h0;
      else \nr00071[1] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [4] <= 1'h0;
      else \nr00071[1] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [5] <= 1'h0;
      else \nr00071[1] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [6] <= 1'h0;
      else \nr00071[1] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [7] <= 1'h0;
      else \nr00071[1] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [8] <= 1'h0;
      else \nr00071[1] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [9] <= 1'h0;
      else \nr00071[1] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [10] <= 1'h0;
      else \nr00071[1] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [11] <= 1'h0;
      else \nr00071[1] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [12] <= 1'h0;
      else \nr00071[1] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [13] <= 1'h0;
      else \nr00071[1] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [14] <= 1'h0;
      else \nr00071[1] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [15] <= 1'h0;
      else \nr00071[1] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [16] <= 1'h0;
      else \nr00071[1] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [17] <= 1'h0;
      else \nr00071[1] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [18] <= 1'h0;
      else \nr00071[1] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [19] <= 1'h0;
      else \nr00071[1] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [20] <= 1'h0;
      else \nr00071[1] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [21] <= 1'h0;
      else \nr00071[1] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [22] <= 1'h0;
      else \nr00071[1] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [23] <= 1'h0;
      else \nr00071[1] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [24] <= 1'h0;
      else \nr00071[1] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [25] <= 1'h0;
      else \nr00071[1] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [26] <= 1'h0;
      else \nr00071[1] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [27] <= 1'h0;
      else \nr00071[1] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [28] <= 1'h0;
      else \nr00071[1] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [29] <= 1'h0;
      else \nr00071[1] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [30] <= 1'h0;
      else \nr00071[1] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00029)
      if (!nw00395) \nr00071[1] [31] <= 1'h0;
      else \nr00071[1] [31] <= nw00089;
  reg \nr00123[0] ;
  always @(posedge clock_10_i)
    \nr00123[0]  <= nw00006;
  assign nw05430[0] = \nr00123[0] ;
  reg \nr00123[1] ;
  always @(posedge clock_10_i)
    \nr00123[1]  <= nw00007;
  assign nw05430[1] = \nr00123[1] ;
  reg \nr00123[2] ;
  always @(posedge clock_10_i)
    \nr00123[2]  <= nw00008;
  assign nw05430[2] = \nr00123[2] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00011u  <= nw00052;
  always @(posedge clock_10_i)
    if (nw00041) \nr00011  <= nw00053;
  always @(posedge clock_10_i)
    if (nw00041) \nr00010  <= nw00051;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [0] <= nw00202;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [1] <= nw00213;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [2] <= nw00224;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [3] <= nw00227;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [4] <= nw00228;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [5] <= nw00229;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [6] <= nw00230;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [7] <= nw00231;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [8] <= nw00232;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [9] <= nw00233;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [10] <= nw00203;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [11] <= nw00204;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [12] <= nw00205;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [13] <= nw00206;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [14] <= nw00207;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [15] <= nw00208;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [16] <= nw00209;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [17] <= nw00210;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [18] <= nw00211;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [19] <= nw00212;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [20] <= nw00214;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [21] <= nw00215;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [22] <= nw00216;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [23] <= nw00217;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [24] <= nw00218;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [25] <= nw00219;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [26] <= nw00220;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [27] <= nw00221;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [28] <= nw00222;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [29] <= nw00223;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [30] <= nw00225;
  always @(posedge clock_10_i)
    if (nw00042) \nr00014 [31] <= nw00226;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [0] <= nw00170;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [1] <= nw00181;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [2] <= nw00192;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [3] <= nw00195;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [4] <= nw00196;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [5] <= nw00197;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [6] <= nw00198;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [7] <= nw00199;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [8] <= nw00200;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [9] <= nw00201;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [10] <= nw00171;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [11] <= nw00172;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [12] <= nw00173;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [13] <= nw00174;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [14] <= nw00175;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [15] <= nw00176;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [16] <= nw00177;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [17] <= nw00178;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [18] <= nw00179;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [19] <= nw00180;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [20] <= nw00182;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [21] <= nw00183;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [22] <= nw00184;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [23] <= nw00185;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [24] <= nw00186;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [25] <= nw00187;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [26] <= nw00188;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [27] <= nw00189;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [28] <= nw00190;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [29] <= nw00191;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [30] <= nw00193;
  always @(posedge clock_10_i)
    if (nw00042) \nr00013 [31] <= nw00194;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [0] <= nw00317;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [1] <= nw00328;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [2] <= nw00339;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [3] <= nw00342;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [4] <= nw00343;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [5] <= nw00344;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [6] <= nw00345;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [7] <= nw00346;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [8] <= nw00347;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [9] <= nw00348;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [10] <= nw00318;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [11] <= nw00319;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [12] <= nw00320;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [13] <= nw00321;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [14] <= nw00322;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [15] <= nw00323;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [16] <= nw00324;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [17] <= nw00325;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [18] <= nw00326;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [19] <= nw00327;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [20] <= nw00329;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [21] <= nw00330;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [22] <= nw00331;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [23] <= nw00332;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [24] <= nw00333;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [25] <= nw00334;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [26] <= nw00335;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [27] <= nw00336;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [28] <= nw00337;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [29] <= nw00338;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [30] <= nw00340;
  always @(posedge clock_10_i)
    if (nw00042) \nr00016 [31] <= nw00341;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [5] <= 1'h0;
      else \nr00017 [5] <= nw00312;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [6] <= 1'h0;
      else \nr00017 [6] <= nw00313;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [7] <= 1'h0;
      else \nr00017 [7] <= nw00314;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [8] <= 1'h0;
      else \nr00017 [8] <= nw00315;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [9] <= 1'h0;
      else \nr00017 [9] <= nw00316;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [10] <= 1'h0;
      else \nr00017 [10] <= nw00290;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [11] <= 1'h0;
      else \nr00017 [11] <= nw00291;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [12] <= 1'h0;
      else \nr00017 [12] <= nw00292;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [13] <= 1'h0;
      else \nr00017 [13] <= nw00293;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [14] <= 1'h0;
      else \nr00017 [14] <= nw00294;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [15] <= 1'h0;
      else \nr00017 [15] <= nw00295;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [16] <= 1'h0;
      else \nr00017 [16] <= nw00296;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [17] <= 1'h0;
      else \nr00017 [17] <= nw00297;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [18] <= 1'h0;
      else \nr00017 [18] <= nw00298;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [19] <= 1'h0;
      else \nr00017 [19] <= nw00299;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [20] <= 1'h0;
      else \nr00017 [20] <= nw00300;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [21] <= 1'h0;
      else \nr00017 [21] <= nw00301;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [22] <= 1'h0;
      else \nr00017 [22] <= nw00302;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [23] <= 1'h0;
      else \nr00017 [23] <= nw00303;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [24] <= 1'h0;
      else \nr00017 [24] <= nw00304;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [25] <= 1'h0;
      else \nr00017 [25] <= nw00305;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [26] <= 1'h0;
      else \nr00017 [26] <= nw00306;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [27] <= 1'h0;
      else \nr00017 [27] <= nw00307;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [28] <= 1'h0;
      else \nr00017 [28] <= nw00308;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [29] <= 1'h0;
      else \nr00017 [29] <= nw00309;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [30] <= 1'h0;
      else \nr00017 [30] <= nw00310;
  always @(posedge clock_10_i)
    if (nw00042)
      if (\nw05426 ) \nr00017 [31] <= 1'h0;
      else \nr00017 [31] <= nw00311;
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [1] <= nw05412[1];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [2] <= nw05412[2];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [3] <= nw05412[3];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [4] <= nw05412[4];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [5] <= nw05412[5];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [6] <= nw05412[6];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [7] <= nw05412[7];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [8] <= nw05412[8];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [9] <= nw05412[9];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [10] <= nw05412[10];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [11] <= nw05412[11];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [12] <= nw05412[12];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [13] <= nw05412[13];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [14] <= nw05412[14];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [15] <= nw05412[15];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [16] <= nw05412[16];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [17] <= nw05412[17];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [18] <= nw05412[18];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [19] <= nw05412[19];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [20] <= nw05412[20];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [21] <= nw05412[21];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [22] <= nw05412[22];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [23] <= nw05412[23];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [24] <= nw05412[24];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [25] <= nw05412[25];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [26] <= nw05412[26];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [27] <= nw05412[27];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [28] <= nw05412[28];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [29] <= nw05412[29];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [30] <= nw05412[30];
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [31] <= nw05412[31];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [0] <= nw05409[0];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [1] <= nw05409[1];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [2] <= nw05409[2];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [3] <= nw05409[3];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [4] <= nw05409[4];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [5] <= nw05409[5];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [6] <= nw05409[6];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [7] <= nw05409[7];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [8] <= nw05409[8];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [9] <= nw05409[9];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [10] <= nw05409[10];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [11] <= nw05409[11];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [12] <= nw05409[12];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [13] <= nw05409[13];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [14] <= nw05409[14];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [15] <= nw05409[15];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [16] <= nw05409[16];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [17] <= nw05409[17];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [18] <= nw05409[18];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [19] <= nw05409[19];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [20] <= nw05409[20];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [21] <= nw05409[21];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [22] <= nw05409[22];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [23] <= nw05409[23];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [24] <= nw05409[24];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [25] <= nw05409[25];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [26] <= nw05409[26];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [27] <= nw05409[27];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [28] <= nw05409[28];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [29] <= nw05409[29];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [30] <= nw05409[30];
  always @(posedge clock_10_i)
    if (nw00041) \nr00024 [31] <= nw05409[31];
  reg \nr00126[0] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[0]  <= nw05419[0];
  assign \nw05422 [0] = \nr00126[0] ;
  reg \nr00126[1] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[1]  <= nw05419[1];
  assign \nw05422 [1] = \nr00126[1] ;
  reg \nr00126[2] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[2]  <= nw05419[2];
  assign \nw05422 [2] = \nr00126[2] ;
  reg \nr00126[3] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[3]  <= nw05419[3];
  assign \nw05422 [3] = \nr00126[3] ;
  reg \nr00126[4] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[4]  <= nw05419[4];
  assign \nw05422 [4] = \nr00126[4] ;
  reg \nr00126[5] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[5]  <= nw05419[5];
  assign \nw05422 [5] = \nr00126[5] ;
  reg \nr00126[6] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[6]  <= nw05419[6];
  assign \nw05422 [6] = \nr00126[6] ;
  reg \nr00126[7] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[7]  <= nw05419[7];
  assign \nw05422 [7] = \nr00126[7] ;
  reg \nr00126[8] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[8]  <= nw05419[8];
  assign \nw05422 [8] = \nr00126[8] ;
  reg \nr00126[9] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[9]  <= nw05419[9];
  assign \nw05422 [9] = \nr00126[9] ;
  reg \nr00126[10] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[10]  <= nw05419[10];
  assign \nw05422 [10] = \nr00126[10] ;
  reg \nr00126[11] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[11]  <= nw05419[11];
  assign \nw05422 [11] = \nr00126[11] ;
  reg \nr00126[12] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[12]  <= nw05419[12];
  assign \nw05422 [12] = \nr00126[12] ;
  reg \nr00126[13] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[13]  <= nw05419[13];
  assign \nw05422 [13] = \nr00126[13] ;
  reg \nr00126[14] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[14]  <= nw05419[14];
  assign \nw05422 [14] = \nr00126[14] ;
  reg \nr00126[15] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[15]  <= nw05419[15];
  assign \nw05422 [15] = \nr00126[15] ;
  reg \nr00126[16] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[16]  <= nw05419[16];
  assign \nw05422 [16] = \nr00126[16] ;
  reg \nr00126[17] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[17]  <= nw05419[17];
  assign \nw05422 [17] = \nr00126[17] ;
  reg \nr00126[18] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[18]  <= nw05419[18];
  assign \nw05422 [18] = \nr00126[18] ;
  reg \nr00126[19] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[19]  <= nw05419[19];
  assign \nw05422 [19] = \nr00126[19] ;
  reg \nr00126[20] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[20]  <= nw05419[20];
  assign \nw05422 [20] = \nr00126[20] ;
  reg \nr00126[21] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[21]  <= nw05419[21];
  assign \nw05422 [21] = \nr00126[21] ;
  reg \nr00126[22] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[22]  <= nw05419[22];
  assign \nw05422 [22] = \nr00126[22] ;
  reg \nr00126[23] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[23]  <= nw05419[23];
  assign \nw05422 [23] = \nr00126[23] ;
  reg \nr00126[24] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[24]  <= nw05419[24];
  assign \nw05422 [24] = \nr00126[24] ;
  reg \nr00126[25] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[25]  <= nw05419[25];
  assign \nw05422 [25] = \nr00126[25] ;
  reg \nr00126[26] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[26]  <= nw05419[26];
  assign \nw05422 [26] = \nr00126[26] ;
  reg \nr00126[27] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[27]  <= nw05419[27];
  assign \nw05422 [27] = \nr00126[27] ;
  reg \nr00126[28] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[28]  <= nw05419[28];
  assign \nw05422 [28] = \nr00126[28] ;
  reg \nr00126[29] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[29]  <= nw05419[29];
  assign \nw05422 [29] = \nr00126[29] ;
  reg \nr00126[30] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[30]  <= nw05419[30];
  assign \nw05422 [30] = \nr00126[30] ;
  reg \nr00126[31] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00126[31]  <= nw05419[31];
  assign \nw05422 [31] = \nr00126[31] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [16] <= nw05418[16];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [17] <= nw05418[17];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [18] <= nw05418[18];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [19] <= nw05418[19];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [20] <= nw05418[20];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [21] <= nw05418[21];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [22] <= nw05418[22];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [23] <= nw05418[23];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [24] <= nw05418[24];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [25] <= nw05418[25];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [26] <= nw05418[26];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [27] <= nw05418[27];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [28] <= nw05418[28];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [29] <= nw05418[29];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [30] <= nw05418[30];
  always @(posedge clock_10_i)
    if (nw00041) \nr00021 [31] <= nw05418[31];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [0] <= nw05410[0];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [1] <= nw05413[1];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [2] <= nw05413[2];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [3] <= nw05413[3];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [4] <= nw05413[4];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [5] <= nw05413[5];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [6] <= nw05413[6];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [7] <= nw05413[7];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [8] <= nw05413[8];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [9] <= nw05413[9];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [10] <= nw05413[10];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [11] <= nw05413[11];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [12] <= nw05413[12];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [13] <= nw05413[13];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [14] <= nw05413[14];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [15] <= nw05413[15];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [16] <= nw05413[16];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [17] <= nw05413[17];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [18] <= nw05413[18];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [19] <= nw05413[19];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [20] <= nw05413[20];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [21] <= nw05413[21];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [22] <= nw05413[22];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [23] <= nw05413[23];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [24] <= nw05413[24];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [25] <= nw05413[25];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [26] <= nw05413[26];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [27] <= nw05413[27];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [28] <= nw05413[28];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [29] <= nw05413[29];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [30] <= nw05413[30];
  always @(posedge clock_10_i)
    if (nw00041) \nr00019 [31] <= nw05413[31];
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [0] <= nw00234;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [1] <= nw00245;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [2] <= nw00256;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [3] <= nw00259;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [4] <= nw00260;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [5] <= nw00261;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [6] <= nw00262;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [7] <= nw00263;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [8] <= nw00264;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [9] <= nw00265;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [10] <= nw00235;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [11] <= nw00236;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [12] <= nw00237;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [13] <= nw00238;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [14] <= nw00239;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [15] <= nw00240;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [16] <= nw00241;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [17] <= nw00242;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [18] <= nw00243;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [19] <= nw00244;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [20] <= nw00246;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [21] <= nw00247;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [22] <= nw00248;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [23] <= nw00249;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [24] <= nw00250;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [25] <= nw00251;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [26] <= nw00252;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [27] <= nw00253;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [28] <= nw00254;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [29] <= nw00255;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [30] <= nw00257;
  always @(posedge clock_10_i)
    if (nw00041) \nr00020 [31] <= nw00258;
  always @(posedge clock_10_i)
    if (nw00041) \nr00018 [0] <= nw05411[0];
  reg \nr00158[1] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[1]  <= nw05411[1];
  assign \nw05423 [1] = \nr00158[1] ;
  reg \nr00158[2] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[2]  <= nw05411[2];
  assign \nw05423 [2] = \nr00158[2] ;
  reg \nr00158[3] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[3]  <= nw05411[3];
  assign \nw05423 [3] = \nr00158[3] ;
  reg \nr00158[4] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[4]  <= nw05411[4];
  assign \nw05423 [4] = \nr00158[4] ;
  reg \nr00158[5] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[5]  <= nw05411[5];
  assign \nw05423 [5] = \nr00158[5] ;
  reg \nr00158[6] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[6]  <= nw05411[6];
  assign \nw05423 [6] = \nr00158[6] ;
  reg \nr00158[7] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[7]  <= nw05411[7];
  assign \nw05423 [7] = \nr00158[7] ;
  reg \nr00158[8] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[8]  <= nw05411[8];
  assign \nw05423 [8] = \nr00158[8] ;
  reg \nr00158[9] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[9]  <= nw05411[9];
  assign \nw05423 [9] = \nr00158[9] ;
  reg \nr00158[10] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[10]  <= nw05411[10];
  assign \nw05423 [10] = \nr00158[10] ;
  reg \nr00158[11] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[11]  <= nw05411[11];
  assign \nw05423 [11] = \nr00158[11] ;
  reg \nr00158[12] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[12]  <= nw05411[12];
  assign \nw05423 [12] = \nr00158[12] ;
  reg \nr00158[13] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[13]  <= nw05411[13];
  assign \nw05423 [13] = \nr00158[13] ;
  reg \nr00158[14] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[14]  <= nw05411[14];
  assign \nw05423 [14] = \nr00158[14] ;
  reg \nr00158[15] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[15]  <= nw05411[15];
  assign \nw05423 [15] = \nr00158[15] ;
  reg \nr00158[16] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[16]  <= nw05411[16];
  assign \nw05423 [16] = \nr00158[16] ;
  reg \nr00158[17] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[17]  <= nw05411[17];
  assign \nw05423 [17] = \nr00158[17] ;
  reg \nr00158[18] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[18]  <= nw05411[18];
  assign \nw05423 [18] = \nr00158[18] ;
  reg \nr00158[19] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[19]  <= nw05411[19];
  assign \nw05423 [19] = \nr00158[19] ;
  reg \nr00158[20] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[20]  <= nw05411[20];
  assign \nw05423 [20] = \nr00158[20] ;
  reg \nr00158[21] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[21]  <= nw05411[21];
  assign \nw05423 [21] = \nr00158[21] ;
  reg \nr00158[22] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[22]  <= nw05411[22];
  assign \nw05423 [22] = \nr00158[22] ;
  reg \nr00158[23] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[23]  <= nw05411[23];
  assign \nw05423 [23] = \nr00158[23] ;
  reg \nr00158[24] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[24]  <= nw05411[24];
  assign \nw05423 [24] = \nr00158[24] ;
  reg \nr00158[25] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[25]  <= nw05411[25];
  assign \nw05423 [25] = \nr00158[25] ;
  reg \nr00158[26] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[26]  <= nw05411[26];
  assign \nw05423 [26] = \nr00158[26] ;
  reg \nr00158[27] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[27]  <= nw05411[27];
  assign \nw05423 [27] = \nr00158[27] ;
  reg \nr00158[28] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[28]  <= nw05411[28];
  assign \nw05423 [28] = \nr00158[28] ;
  reg \nr00158[29] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[29]  <= nw05411[29];
  assign \nw05423 [29] = \nr00158[29] ;
  reg \nr00158[30] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[30]  <= nw05411[30];
  assign \nw05423 [30] = \nr00158[30] ;
  reg \nr00158[31] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00158[31]  <= nw05411[31];
  assign \nw05423 [31] = \nr00158[31] ;
  always @(posedge clock_10_i)
    if (nw00041) \nr00021tu  <= nw00050;
  always @(posedge clock_10_i)
    if (nw00041) \nr00021t  <= nw00054;
  always @(posedge clock_10_i)
    if (nw00043) \nr00037  <= nw00137;
  always @(posedge clock_10_i)
    if (nw00043) \nr00060  <= nw00136;
  always @(posedge clock_10_i)
    if (nw00043) \nr00049  <= nw00135;
  always @(posedge clock_10_i)
    if (nw00043) \nr00048  <= nw00134;
  always @(posedge clock_10_i)
    if (nw00043) \nr00042U  <= nw00133;
  always @(posedge clock_10_i)
    if (nw00043) \nr00040U  <= nw00132;
  always @(posedge clock_10_i)
    if (nw00043) \nr00045  <= nw00131;
  always @(posedge clock_10_i)
    if (nw00043) \nr00042  <= nw00130;
  always @(posedge clock_10_i)
    if (nw00043) \nr00040  <= nw00129;
  always @(posedge clock_10_i)
    if (nw00043) \nr00028  <= nw00128;
  always @(posedge clock_10_i)
    if (nw00043) \nr00046  <= nw00127;
  always @(posedge clock_10_i)
    if (nw00043) \nr00056  <= nw00126;
  always @(posedge clock_10_i)
    if (nw00043) \nr00058  <= nw00125;
  always @(posedge clock_10_i)
    if (nw00043) \nr00061  <= nw00124;
  always @(posedge clock_10_i)
    if (nw00043) \nr00052U  <= nw00123;
  always @(posedge clock_10_i)
    if (nw00043) \nr00052  <= nw00122;
  always @(posedge clock_10_i)
    if (nw00043) \nr00050  <= nw00121;
  always @(posedge clock_10_i)
    if (nw00043) \nr00015  <= nw00120;
  always @(posedge clock_10_i)
    if (nw00043) \nr00027  <= nw00119;
  always @(posedge clock_10_i)
    if (nw00043) \nr00056I  <= nw00118;
  always @(posedge clock_10_i)
    if (nw00043) \nr00058I  <= nw00117;
  always @(posedge clock_10_i)
    if (nw00043) \nr00050I  <= nw00116;
  always @(posedge clock_10_i)
    if (nw00043) \nr00028I  <= nw00115;
  always @(posedge clock_10_i)
    if (nw00043) \nr00046I  <= nw00114;
  always @(posedge clock_10_i)
    if (nw00043) \nr00061I  <= nw00113;
  always @(posedge clock_10_i)
    if (nw00043) \nr00052IU  <= nw00112;
  always @(posedge clock_10_i)
    if (nw00043) \nr00052I  <= nw00111;
  always @(posedge clock_10_i)
    if (nw00043) \nr00032U  <= nw00110;
  always @(posedge clock_10_i)
    if (nw00043) \nr00034U  <= nw00109;
  always @(posedge clock_10_i)
    if (nw00043) \nr00032  <= nw00108;
  always @(posedge clock_10_i)
    if (nw00043) \nr00034  <= nw00107;
  always @(posedge clock_10_i)
    if (nw00043) \nr00036  <= nw00106;
  always @(posedge clock_10_i)
    if (nw00043) \nr00031  <= nw00105;
  always @(posedge clock_10_i)
    if (nw00043) \nr00038R  <= nw00104;
  always @(posedge clock_10_i)
    if (nw00043) \nr00038  <= nw05416[0];
  always @(posedge clock_10_i)
    if (nw00043) \nr00030  <= nw00103;
  always @(posedge clock_10_i)
    if (nw00043) \nr00044  <= nw00102;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00063  <= 1'h0;
    else \nr00063  <= nw00349;
  always @(posedge clock_10_i)
    if (\nw05425 ) nr00008 <= 1'h0;
    else nr00008 <= nw00350;
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [0] <= \nw05424 [0];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [1] <= \nw05424 [1];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [2] <= \nw05424 [2];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [3] <= \nw05424 [3];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [4] <= \nw05424 [4];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [5] <= \nw05424 [5];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [6] <= \nw05424 [6];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [7] <= \nw05424 [7];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [8] <= \nw05424 [8];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [9] <= \nw05424 [9];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [10] <= \nw05424 [10];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [11] <= \nw05424 [11];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [12] <= \nw05424 [12];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [13] <= \nw05424 [13];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [14] <= \nw05424 [14];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [15] <= \nw05424 [15];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [16] <= \nw05424 [16];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [17] <= \nw05424 [17];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [18] <= \nw05424 [18];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [19] <= \nw05424 [19];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [20] <= \nw05424 [20];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [21] <= \nw05424 [21];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [22] <= \nw05424 [22];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [23] <= \nw05424 [23];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [24] <= \nw05424 [24];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [25] <= \nw05424 [25];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [26] <= \nw05424 [26];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [27] <= \nw05424 [27];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [28] <= \nw05424 [28];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [29] <= \nw05424 [29];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [30] <= \nw05424 [30];
  always @(posedge clock_10_i)
    if (nw00045) \nr00064 [31] <= \nw05424 [31];
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[0] <= 1'h0;
    else if (nw00044) ext_bus_data_o[0] <= nw00202;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[1] <= 1'h0;
    else if (nw00044) ext_bus_data_o[1] <= nw00213;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[2] <= 1'h0;
    else if (nw00044) ext_bus_data_o[2] <= nw00224;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[3] <= 1'h0;
    else if (nw00044) ext_bus_data_o[3] <= nw00227;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[4] <= 1'h0;
    else if (nw00044) ext_bus_data_o[4] <= nw00228;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[5] <= 1'h0;
    else if (nw00044) ext_bus_data_o[5] <= nw00229;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[6] <= 1'h0;
    else if (nw00044) ext_bus_data_o[6] <= nw00230;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[7] <= 1'h0;
    else if (nw00044) ext_bus_data_o[7] <= nw00231;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[8] <= 1'h0;
    else if (nw00044) ext_bus_data_o[8] <= nw00274;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[9] <= 1'h0;
    else if (nw00044) ext_bus_data_o[9] <= nw00275;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[10] <= 1'h0;
    else if (nw00044) ext_bus_data_o[10] <= nw00276;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[11] <= 1'h0;
    else if (nw00044) ext_bus_data_o[11] <= nw00277;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[12] <= 1'h0;
    else if (nw00044) ext_bus_data_o[12] <= nw00278;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[13] <= 1'h0;
    else if (nw00044) ext_bus_data_o[13] <= nw00279;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[14] <= 1'h0;
    else if (nw00044) ext_bus_data_o[14] <= nw00280;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[15] <= 1'h0;
    else if (nw00044) ext_bus_data_o[15] <= nw00281;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[16] <= 1'h0;
    else if (nw00044) ext_bus_data_o[16] <= nw00282;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[17] <= 1'h0;
    else if (nw00044) ext_bus_data_o[17] <= nw00283;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[18] <= 1'h0;
    else if (nw00044) ext_bus_data_o[18] <= nw00284;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[19] <= 1'h0;
    else if (nw00044) ext_bus_data_o[19] <= nw00285;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[20] <= 1'h0;
    else if (nw00044) ext_bus_data_o[20] <= nw00286;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[21] <= 1'h0;
    else if (nw00044) ext_bus_data_o[21] <= nw00287;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[22] <= 1'h0;
    else if (nw00044) ext_bus_data_o[22] <= nw00288;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[23] <= 1'h0;
    else if (nw00044) ext_bus_data_o[23] <= nw00289;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[24] <= 1'h0;
    else if (nw00044) ext_bus_data_o[24] <= nw00266;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[25] <= 1'h0;
    else if (nw00044) ext_bus_data_o[25] <= nw00267;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[26] <= 1'h0;
    else if (nw00044) ext_bus_data_o[26] <= nw00268;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[27] <= 1'h0;
    else if (nw00044) ext_bus_data_o[27] <= nw00269;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[28] <= 1'h0;
    else if (nw00044) ext_bus_data_o[28] <= nw00270;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[29] <= 1'h0;
    else if (nw00044) ext_bus_data_o[29] <= nw00271;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[30] <= 1'h0;
    else if (nw00044) ext_bus_data_o[30] <= nw00272;
  always @(posedge clock_10_i)
    if (\nw05425 ) ext_bus_data_o[31] <= 1'h0;
    else if (nw00044) ext_bus_data_o[31] <= nw00273;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00065  <= 1'h0;
    else \nr00065  <= nw00383;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[0] <= 1'h0;
    else if (nw00046) address_ext_o[0] <= nw00351;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[1] <= 1'h0;
    else if (nw00046) address_ext_o[1] <= nw00362;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[2] <= 1'h0;
    else if (nw00046) address_ext_o[2] <= nw00373;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[3] <= 1'h0;
    else if (nw00046) address_ext_o[3] <= nw00376;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[4] <= 1'h0;
    else if (nw00046) address_ext_o[4] <= nw00377;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[5] <= 1'h0;
    else if (nw00046) address_ext_o[5] <= nw00378;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[6] <= 1'h0;
    else if (nw00046) address_ext_o[6] <= nw00379;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[7] <= 1'h0;
    else if (nw00046) address_ext_o[7] <= nw00380;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[8] <= 1'h0;
    else if (nw00046) address_ext_o[8] <= nw00381;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[9] <= 1'h0;
    else if (nw00046) address_ext_o[9] <= nw00382;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[10] <= 1'h0;
    else if (nw00046) address_ext_o[10] <= nw00352;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[11] <= 1'h0;
    else if (nw00046) address_ext_o[11] <= nw00353;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[12] <= 1'h0;
    else if (nw00046) address_ext_o[12] <= nw00354;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[13] <= 1'h0;
    else if (nw00046) address_ext_o[13] <= nw00355;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[14] <= 1'h0;
    else if (nw00046) address_ext_o[14] <= nw00356;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[15] <= 1'h0;
    else if (nw00046) address_ext_o[15] <= nw00357;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[16] <= 1'h0;
    else if (nw00046) address_ext_o[16] <= nw00358;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[17] <= 1'h0;
    else if (nw00046) address_ext_o[17] <= nw00359;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[18] <= 1'h0;
    else if (nw00046) address_ext_o[18] <= nw00360;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[19] <= 1'h0;
    else if (nw00046) address_ext_o[19] <= nw00361;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[20] <= 1'h0;
    else if (nw00046) address_ext_o[20] <= nw00363;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[21] <= 1'h0;
    else if (nw00046) address_ext_o[21] <= nw00364;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[22] <= 1'h0;
    else if (nw00046) address_ext_o[22] <= nw00365;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[23] <= 1'h0;
    else if (nw00046) address_ext_o[23] <= nw00366;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[24] <= 1'h0;
    else if (nw00046) address_ext_o[24] <= nw00367;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[25] <= 1'h0;
    else if (nw00046) address_ext_o[25] <= nw00368;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[26] <= 1'h0;
    else if (nw00046) address_ext_o[26] <= nw00369;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[27] <= 1'h0;
    else if (nw00046) address_ext_o[27] <= nw00370;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[28] <= 1'h0;
    else if (nw00046) address_ext_o[28] <= nw00371;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[29] <= 1'h0;
    else if (nw00046) address_ext_o[29] <= nw00372;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[30] <= 1'h0;
    else if (nw00046) address_ext_o[30] <= nw00374;
  always @(posedge clock_10_i)
    if (\nw05425 ) address_ext_o[31] <= 1'h0;
    else if (nw00046) address_ext_o[31] <= nw00375;
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [0] <= nw05417[0];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [1] <= nw05417[1];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [2] <= nw05417[2];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [3] <= nw05417[3];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [4] <= nw05417[4];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [5] <= nw05417[5];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [6] <= nw05417[6];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [7] <= nw05417[7];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [8] <= nw05417[8];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [9] <= nw05417[9];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [10] <= nw05417[10];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [11] <= nw05417[11];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [12] <= nw05417[12];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [13] <= nw05417[13];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [14] <= nw05417[14];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [15] <= nw05417[15];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [16] <= nw05417[16];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [17] <= nw05417[17];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [18] <= nw05417[18];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [19] <= nw05417[19];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [20] <= nw05417[20];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [21] <= nw05417[21];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [22] <= nw05417[22];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [23] <= nw05417[23];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [24] <= nw05417[24];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [25] <= nw05417[25];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [26] <= nw05417[26];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [27] <= nw05417[27];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [28] <= nw05417[28];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [29] <= nw05417[29];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [30] <= nw05417[30];
  always @(posedge clock_10_i)
    if (nw00043) \nr00026 [31] <= \nr00064 [31];
  always @(posedge clock_10_i)
    if (nw00043) \nr00068 [0] <= \nr00064 [7];
  always @(posedge clock_10_i)
    if (nw00043) \nr00068 [1] <= \nr00064 [8];
  always @(posedge clock_10_i)
    if (nw00043) \nr00068 [2] <= \nr00064 [9];
  always @(posedge clock_10_i)
    if (nw00043) \nr00068 [3] <= \nr00064 [10];
  always @(posedge clock_10_i)
    if (nw00043) \nr00068 [4] <= \nr00064 [11];
  always @(posedge clock_10_i)
    if (nw00043) \nr00070 [0] <= \nr00064 [20];
  always @(posedge clock_10_i)
    if (nw00043) \nr00070 [1] <= \nr00064 [21];
  always @(posedge clock_10_i)
    if (nw00043) \nr00070 [2] <= \nr00064 [22];
  always @(posedge clock_10_i)
    if (nw00043) \nr00070 [3] <= \nr00064 [23];
  always @(posedge clock_10_i)
    if (nw00043) \nr00070 [4] <= \nr00064 [24];
  always @(posedge clock_10_i)
    if (nw00043) \nr00069 [0] <= \nr00064 [15];
  always @(posedge clock_10_i)
    if (nw00043) \nr00069 [1] <= \nr00064 [16];
  always @(posedge clock_10_i)
    if (nw00043) \nr00069 [2] <= \nr00064 [17];
  always @(posedge clock_10_i)
    if (nw00043) \nr00069 [3] <= \nr00064 [18];
  always @(posedge clock_10_i)
    if (nw00043) \nr00069 [4] <= \nr00064 [19];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [0] <= 1'h0;
    else if (nw00048) \nr00067 [0] <= \nr00066 [0];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [1] <= 1'h0;
    else if (nw00048) \nr00067 [1] <= \nr00066 [1];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [2] <= 1'h0;
    else if (nw00048) \nr00067 [2] <= \nr00066 [2];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [3] <= 1'h0;
    else if (nw00048) \nr00067 [3] <= \nr00066 [3];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [4] <= 1'h0;
    else if (nw00048) \nr00067 [4] <= \nr00066 [4];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [5] <= 1'h0;
    else if (nw00048) \nr00067 [5] <= \nr00066 [5];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [6] <= 1'h0;
    else if (nw00048) \nr00067 [6] <= \nr00066 [6];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [7] <= 1'h0;
    else if (nw00048) \nr00067 [7] <= \nr00066 [7];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [8] <= 1'h0;
    else if (nw00048) \nr00067 [8] <= \nr00066 [8];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [9] <= 1'h0;
    else if (nw00048) \nr00067 [9] <= \nr00066 [9];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [10] <= 1'h0;
    else if (nw00048) \nr00067 [10] <= \nr00066 [10];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [11] <= 1'h0;
    else if (nw00048) \nr00067 [11] <= \nr00066 [11];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [12] <= 1'h0;
    else if (nw00048) \nr00067 [12] <= \nr00066 [12];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [13] <= 1'h0;
    else if (nw00048) \nr00067 [13] <= \nr00066 [13];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [14] <= 1'h0;
    else if (nw00048) \nr00067 [14] <= \nr00066 [14];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [15] <= 1'h0;
    else if (nw00048) \nr00067 [15] <= \nr00066 [15];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [16] <= 1'h0;
    else if (nw00048) \nr00067 [16] <= \nr00066 [16];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [17] <= 1'h0;
    else if (nw00048) \nr00067 [17] <= \nr00066 [17];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [18] <= 1'h0;
    else if (nw00048) \nr00067 [18] <= \nr00066 [18];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [19] <= 1'h0;
    else if (nw00048) \nr00067 [19] <= \nr00066 [19];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [20] <= 1'h0;
    else if (nw00048) \nr00067 [20] <= \nr00066 [20];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [21] <= 1'h0;
    else if (nw00048) \nr00067 [21] <= \nr00066 [21];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [22] <= 1'h0;
    else if (nw00048) \nr00067 [22] <= \nr00066 [22];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [23] <= 1'h0;
    else if (nw00048) \nr00067 [23] <= \nr00066 [23];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [24] <= 1'h0;
    else if (nw00048) \nr00067 [24] <= \nr00066 [24];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [25] <= 1'h0;
    else if (nw00048) \nr00067 [25] <= \nr00066 [25];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [26] <= 1'h0;
    else if (nw00048) \nr00067 [26] <= \nr00066 [26];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [27] <= 1'h0;
    else if (nw00048) \nr00067 [27] <= \nr00066 [27];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [28] <= 1'h0;
    else if (nw00048) \nr00067 [28] <= \nr00066 [28];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [29] <= 1'h0;
    else if (nw00048) \nr00067 [29] <= \nr00066 [29];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [30] <= 1'h0;
    else if (nw00048) \nr00067 [30] <= \nr00066 [30];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00067 [31] <= 1'h0;
    else if (nw00048) \nr00067 [31] <= \nr00066 [31];
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [0] <= 1'h0;
    else if (nw00049) \nr00066 [0] <= nw00138;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [1] <= 1'h0;
    else if (nw00049) \nr00066 [1] <= nw00149;
  always @(posedge clock_10_i)
    nr00001[0] <= nw00060;
  always @(posedge clock_10_i)
    nr00001[1] <= nw00061;
  always @(posedge clock_10_i)
    nr00001[2] <= nw00062;
  always @(posedge clock_10_i)
    nr00001[3] <= nw00063;
  always @(posedge clock_10_i)
    nr00001[4] <= nw00064;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [0] <= 1'h0;
      else \nr00071[10] [0] <= nw00065;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [1] <= 1'h0;
      else \nr00071[10] [1] <= nw00076;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [2] <= 1'h0;
      else \nr00071[10] [2] <= nw00087;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [3] <= 1'h0;
      else \nr00071[10] [3] <= nw00090;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [4] <= 1'h0;
      else \nr00071[10] [4] <= nw00091;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [5] <= 1'h0;
      else \nr00071[10] [5] <= nw00092;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [6] <= 1'h0;
      else \nr00071[10] [6] <= nw00093;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [7] <= 1'h0;
      else \nr00071[10] [7] <= nw00094;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [8] <= 1'h0;
      else \nr00071[10] [8] <= nw00095;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [9] <= 1'h0;
      else \nr00071[10] [9] <= nw00096;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [10] <= 1'h0;
      else \nr00071[10] [10] <= nw00066;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [11] <= 1'h0;
      else \nr00071[10] [11] <= nw00067;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [12] <= 1'h0;
      else \nr00071[10] [12] <= nw00068;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [13] <= 1'h0;
      else \nr00071[10] [13] <= nw00069;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [14] <= 1'h0;
      else \nr00071[10] [14] <= nw00070;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [15] <= 1'h0;
      else \nr00071[10] [15] <= nw00071;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [16] <= 1'h0;
      else \nr00071[10] [16] <= nw00072;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [17] <= 1'h0;
      else \nr00071[10] [17] <= nw00073;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [18] <= 1'h0;
      else \nr00071[10] [18] <= nw00074;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [19] <= 1'h0;
      else \nr00071[10] [19] <= nw00075;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [20] <= 1'h0;
      else \nr00071[10] [20] <= nw00077;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [21] <= 1'h0;
      else \nr00071[10] [21] <= nw00078;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [22] <= 1'h0;
      else \nr00071[10] [22] <= nw00079;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [23] <= 1'h0;
      else \nr00071[10] [23] <= nw00080;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [24] <= 1'h0;
      else \nr00071[10] [24] <= nw00081;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [25] <= 1'h0;
      else \nr00071[10] [25] <= nw00082;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [26] <= 1'h0;
      else \nr00071[10] [26] <= nw00083;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [27] <= 1'h0;
      else \nr00071[10] [27] <= nw00084;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [28] <= 1'h0;
      else \nr00071[10] [28] <= nw00085;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [29] <= 1'h0;
      else \nr00071[10] [29] <= nw00086;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [30] <= 1'h0;
      else \nr00071[10] [30] <= nw00088;
  always @(posedge clock_10_i)
    if (nw00039)
      if (!nw00385) \nr00071[10] [31] <= 1'h0;
      else \nr00071[10] [31] <= nw00089;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [2] <= 1'h0;
    else if (nw00047) \nr00066 [2] <= nw00160;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [3] <= 1'h0;
    else if (nw00047) \nr00066 [3] <= nw00163;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [4] <= 1'h0;
    else if (nw00047) \nr00066 [4] <= nw00164;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [5] <= 1'h0;
    else if (nw00047) \nr00066 [5] <= nw00165;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [6] <= 1'h0;
    else if (nw00047) \nr00066 [6] <= nw00166;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [7] <= 1'h0;
    else if (nw00047) \nr00066 [7] <= nw00167;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [8] <= 1'h0;
    else if (nw00047) \nr00066 [8] <= nw00168;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [9] <= 1'h0;
    else if (nw00047) \nr00066 [9] <= nw00169;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [10] <= 1'h0;
    else if (nw00047) \nr00066 [10] <= nw00139;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [11] <= 1'h0;
    else if (nw00047) \nr00066 [11] <= nw00140;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [12] <= 1'h0;
    else if (nw00047) \nr00066 [12] <= nw00141;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [13] <= 1'h0;
    else if (nw00047) \nr00066 [13] <= nw00142;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [14] <= 1'h0;
    else if (nw00047) \nr00066 [14] <= nw00143;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [15] <= 1'h0;
    else if (nw00047) \nr00066 [15] <= nw00144;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [16] <= 1'h0;
    else if (nw00047) \nr00066 [16] <= nw00145;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [17] <= 1'h0;
    else if (nw00047) \nr00066 [17] <= nw00146;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [18] <= 1'h0;
    else if (nw00047) \nr00066 [18] <= nw00147;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [19] <= 1'h0;
    else if (nw00047) \nr00066 [19] <= nw00148;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [20] <= 1'h0;
    else if (nw00047) \nr00066 [20] <= nw00150;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [21] <= 1'h0;
    else if (nw00047) \nr00066 [21] <= nw00151;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [22] <= 1'h0;
    else if (nw00047) \nr00066 [22] <= nw00152;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [23] <= 1'h0;
    else if (nw00047) \nr00066 [23] <= nw00153;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [24] <= 1'h0;
    else if (nw00047) \nr00066 [24] <= nw00154;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [25] <= 1'h0;
    else if (nw00047) \nr00066 [25] <= nw00155;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [26] <= 1'h0;
    else if (nw00047) \nr00066 [26] <= nw00156;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [27] <= 1'h0;
    else if (nw00047) \nr00066 [27] <= nw00157;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [28] <= 1'h0;
    else if (nw00047) \nr00066 [28] <= nw00158;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [29] <= 1'h0;
    else if (nw00047) \nr00066 [29] <= nw00159;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [30] <= 1'h0;
    else if (nw00047) \nr00066 [30] <= nw00161;
  always @(posedge clock_10_i)
    if (\nw05425 ) \nr00066 [31] <= 1'h0;
    else if (nw00047) \nr00066 [31] <= nw00162;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [0] <= 1'h0;
      else \nr00021 [0] <= nw05393;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [1] <= 1'h0;
      else \nr00021 [1] <= nw05394;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [2] <= 1'h0;
      else \nr00021 [2] <= nw05395;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [3] <= 1'h0;
      else \nr00021 [3] <= nw05396;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [4] <= 1'h0;
      else \nr00021 [4] <= nw05397;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [5] <= 1'h0;
      else \nr00021 [5] <= nw05398;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [6] <= 1'h0;
      else \nr00021 [6] <= nw05399;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [7] <= 1'h0;
      else \nr00021 [7] <= nw05400;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [8] <= 1'h0;
      else \nr00021 [8] <= nw05401;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [9] <= 1'h0;
      else \nr00021 [9] <= nw05402;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [10] <= 1'h0;
      else \nr00021 [10] <= nw05403;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [11] <= 1'h0;
      else \nr00021 [11] <= nw05404;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [12] <= 1'h0;
      else \nr00021 [12] <= nw05405;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [13] <= 1'h0;
      else \nr00021 [13] <= nw05406;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [14] <= 1'h0;
      else \nr00021 [14] <= nw05407;
  always @(posedge clock_10_i)
    if (nw00041)
      if (\nr00017 [4]) \nr00021 [15] <= 1'h0;
      else \nr00021 [15] <= nw05408;
  assign nw05412[0] = nw05411[0];
  assign nw05413[0] = nw05410[0];
  assign nw05414[19:1] = \nw05427 [19:1];
  assign nw05415[0] = nw05414[0];
  assign \nw05422 [32] = 1'hx;
  assign \nw05423 [0] = \nr00018 [0];
  assign dp_o = 1'h1;
  assign instr_addr_bus_o = address_ext_o[10:0];
  assign ram_address_bus_o = address_ext_o[9:0];
  assign ram_data_in_o = ext_bus_data_o;
endmodule
